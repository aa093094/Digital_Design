function signed [7:0] conv_kernel;
    input [2:0] i, j;    
    begin
    case({i,j})
     6'b000000: conv_kernel = 8'hdf;
     6'b000001: conv_kernel = 8'hfd;
     6'b000010: conv_kernel = 8'ha;
     6'b000011: conv_kernel = 8'h19;
     6'b000100: conv_kernel = 8'hf6;
     6'b001000: conv_kernel = 8'he6;
     6'b001001: conv_kernel = 8'h1d;
     6'b001010: conv_kernel = 8'h2f;
     6'b001011: conv_kernel = 8'h1a;
     6'b001100: conv_kernel = 8'hd5;
     6'b010000: conv_kernel = 8'h3;
     6'b010001: conv_kernel = 8'h3d;
     6'b010010: conv_kernel = 8'h47;
     6'b010011: conv_kernel = 8'h33;
     6'b010100: conv_kernel = 8'hf2;
     6'b011000: conv_kernel = 8'h17;
     6'b011001: conv_kernel = 8'h12;
     6'b011010: conv_kernel = 8'h2c;
     6'b011011: conv_kernel = 8'h1f;
     6'b011100: conv_kernel = 8'h7;
     6'b100000: conv_kernel = 8'hd3;
     6'b100001: conv_kernel = 8'hcb;
     6'b100010: conv_kernel = 8'hca;
     6'b100011: conv_kernel = 8'hde;
     6'b100100: conv_kernel = 8'he;
     default: conv_kernel = 8'h0;
    endcase
    end
endfunction

function signed [7:0] fc_kernel;
    input [3:0] i;
    input [9:0] j;
    begin
    case({i,j})
     14'b00000000000000: fc_kernel = 8'h06;
     14'b00000000000001: fc_kernel = 8'h01;
     14'b00000000000010: fc_kernel = 8'h05;
     14'b00000000000011: fc_kernel = 8'h04;
     14'b00000000000100: fc_kernel = 8'hf7;
     14'b00000000000101: fc_kernel = 8'h0b;
     14'b00000000000110: fc_kernel = 8'hfe;
     14'b00000000000111: fc_kernel = 8'hf1;
     14'b00000000001000: fc_kernel = 8'hef;
     14'b00000000001001: fc_kernel = 8'h02;
     14'b00000000001010: fc_kernel = 8'h05;
     14'b00000000001011: fc_kernel = 8'h03;
     14'b00000000001100: fc_kernel = 8'hf0;
     14'b00000000001101: fc_kernel = 8'hea;
     14'b00000000001110: fc_kernel = 8'hef;
     14'b00000000001111: fc_kernel = 8'hec;
     14'b00000000010000: fc_kernel = 8'hde;
     14'b00000000010001: fc_kernel = 8'hdf;
     14'b00000000010010: fc_kernel = 8'he4;
     14'b00000000010011: fc_kernel = 8'he1;
     14'b00000000010100: fc_kernel = 8'hf0;
     14'b00000000010101: fc_kernel = 8'hfa;
     14'b00000000010110: fc_kernel = 8'hfd;
     14'b00000000010111: fc_kernel = 8'hf7;
     14'b00000000011000: fc_kernel = 8'h00;
     14'b00000000011001: fc_kernel = 8'h04;
     14'b00000000011010: fc_kernel = 8'h08;
     14'b00000000011011: fc_kernel = 8'he8;
     14'b00000000011100: fc_kernel = 8'hef;
     14'b00000000011101: fc_kernel = 8'hf5;
     14'b00000000011110: fc_kernel = 8'hff;
     14'b00000000011111: fc_kernel = 8'hfc;
     14'b00000000100000: fc_kernel = 8'h00;
     14'b00000000100001: fc_kernel = 8'h03;
     14'b00000000100010: fc_kernel = 8'h00;
     14'b00000000100011: fc_kernel = 8'h05;
     14'b00000000100100: fc_kernel = 8'hfc;
     14'b00000000100101: fc_kernel = 8'h03;
     14'b00000000100110: fc_kernel = 8'hfe;
     14'b00000000100111: fc_kernel = 8'h04;
     14'b00000000101000: fc_kernel = 8'hf9;
     14'b00000000101001: fc_kernel = 8'hfb;
     14'b00000000101010: fc_kernel = 8'hf5;
     14'b00000000101011: fc_kernel = 8'he6;
     14'b00000000101100: fc_kernel = 8'hee;
     14'b00000000101101: fc_kernel = 8'hfc;
     14'b00000000101110: fc_kernel = 8'h06;
     14'b00000000101111: fc_kernel = 8'h01;
     14'b00000000110000: fc_kernel = 8'hf8;
     14'b00000000110001: fc_kernel = 8'h0a;
     14'b00000000110010: fc_kernel = 8'hf1;
     14'b00000000110011: fc_kernel = 8'hd8;
     14'b00000000110100: fc_kernel = 8'hea;
     14'b00000000110101: fc_kernel = 8'hf3;
     14'b00000000110110: fc_kernel = 8'h01;
     14'b00000000110111: fc_kernel = 8'h03;
     14'b00000000111000: fc_kernel = 8'h01;
     14'b00000000111001: fc_kernel = 8'h00;
     14'b00000000111010: fc_kernel = 8'hfa;
     14'b00000000111011: fc_kernel = 8'hfd;
     14'b00000000111100: fc_kernel = 8'hfa;
     14'b00000000111101: fc_kernel = 8'h00;
     14'b00000000111110: fc_kernel = 8'hfc;
     14'b00000000111111: fc_kernel = 8'hfb;
     14'b00000001000000: fc_kernel = 8'hf9;
     14'b00000001000001: fc_kernel = 8'hfb;
     14'b00000001000010: fc_kernel = 8'hf1;
     14'b00000001000011: fc_kernel = 8'hea;
     14'b00000001000100: fc_kernel = 8'he8;
     14'b00000001000101: fc_kernel = 8'hf2;
     14'b00000001000110: fc_kernel = 8'hed;
     14'b00000001000111: fc_kernel = 8'he7;
     14'b00000001001000: fc_kernel = 8'hf0;
     14'b00000001001001: fc_kernel = 8'hf7;
     14'b00000001001010: fc_kernel = 8'hd9;
     14'b00000001001011: fc_kernel = 8'he5;
     14'b00000001001100: fc_kernel = 8'hf5;
     14'b00000001001101: fc_kernel = 8'hff;
     14'b00000001001110: fc_kernel = 8'hfa;
     14'b00000001001111: fc_kernel = 8'hfb;
     14'b00000001010000: fc_kernel = 8'h00;
     14'b00000001010001: fc_kernel = 8'hfd;
     14'b00000001010010: fc_kernel = 8'hfc;
     14'b00000001010011: fc_kernel = 8'hfc;
     14'b00000001010100: fc_kernel = 8'h00;
     14'b00000001010101: fc_kernel = 8'hfe;
     14'b00000001010110: fc_kernel = 8'hfe;
     14'b00000001010111: fc_kernel = 8'h01;
     14'b00000001011000: fc_kernel = 8'h01;
     14'b00000001011001: fc_kernel = 8'hfe;
     14'b00000001011010: fc_kernel = 8'hfb;
     14'b00000001011011: fc_kernel = 8'hff;
     14'b00000001011100: fc_kernel = 8'h00;
     14'b00000001011101: fc_kernel = 8'hf0;
     14'b00000001011110: fc_kernel = 8'he6;
     14'b00000001011111: fc_kernel = 8'hde;
     14'b00000001100000: fc_kernel = 8'hd8;
     14'b00000001100001: fc_kernel = 8'he0;
     14'b00000001100010: fc_kernel = 8'he7;
     14'b00000001100011: fc_kernel = 8'hf4;
     14'b00000001100100: fc_kernel = 8'h01;
     14'b00000001100101: fc_kernel = 8'h02;
     14'b00000001100110: fc_kernel = 8'hf5;
     14'b00000001100111: fc_kernel = 8'hfc;
     14'b00000001101000: fc_kernel = 8'hfd;
     14'b00000001101001: fc_kernel = 8'hfc;
     14'b00000001101010: fc_kernel = 8'hf7;
     14'b00000001101011: fc_kernel = 8'h00;
     14'b00000001101100: fc_kernel = 8'h07;
     14'b00000001101101: fc_kernel = 8'h02;
     14'b00000001101110: fc_kernel = 8'h00;
     14'b00000001101111: fc_kernel = 8'h02;
     14'b00000001110000: fc_kernel = 8'h08;
     14'b00000001110001: fc_kernel = 8'h02;
     14'b00000001110010: fc_kernel = 8'hff;
     14'b00000001110011: fc_kernel = 8'h0a;
     14'b00000001110100: fc_kernel = 8'h04;
     14'b00000001110101: fc_kernel = 8'hf8;
     14'b00000001110110: fc_kernel = 8'he3;
     14'b00000001110111: fc_kernel = 8'hc3;
     14'b00000001111000: fc_kernel = 8'hf6;
     14'b00000001111001: fc_kernel = 8'hd7;
     14'b00000001111010: fc_kernel = 8'hec;
     14'b00000001111011: fc_kernel = 8'hfb;
     14'b00000001111100: fc_kernel = 8'h02;
     14'b00000001111101: fc_kernel = 8'hfe;
     14'b00000001111110: fc_kernel = 8'hf8;
     14'b00000001111111: fc_kernel = 8'hf6;
     14'b00000010000000: fc_kernel = 8'hfe;
     14'b00000010000001: fc_kernel = 8'hfc;
     14'b00000010000010: fc_kernel = 8'h00;
     14'b00000010000011: fc_kernel = 8'h00;
     14'b00000010000100: fc_kernel = 8'h00;
     14'b00000010000101: fc_kernel = 8'hfd;
     14'b00000010000110: fc_kernel = 8'h01;
     14'b00000010000111: fc_kernel = 8'h05;
     14'b00000010001000: fc_kernel = 8'h04;
     14'b00000010001001: fc_kernel = 8'hff;
     14'b00000010001010: fc_kernel = 8'h01;
     14'b00000010001011: fc_kernel = 8'h01;
     14'b00000010001100: fc_kernel = 8'h07;
     14'b00000010001101: fc_kernel = 8'h06;
     14'b00000010001110: fc_kernel = 8'hf1;
     14'b00000010001111: fc_kernel = 8'hc0;
     14'b00000010010000: fc_kernel = 8'h03;
     14'b00000010010001: fc_kernel = 8'hfe;
     14'b00000010010010: fc_kernel = 8'hea;
     14'b00000010010011: fc_kernel = 8'hf9;
     14'b00000010010100: fc_kernel = 8'hfc;
     14'b00000010010101: fc_kernel = 8'hf9;
     14'b00000010010110: fc_kernel = 8'hf6;
     14'b00000010010111: fc_kernel = 8'h03;
     14'b00000010011000: fc_kernel = 8'h02;
     14'b00000010011001: fc_kernel = 8'h00;
     14'b00000010011010: fc_kernel = 8'h03;
     14'b00000010011011: fc_kernel = 8'h01;
     14'b00000010011100: fc_kernel = 8'h01;
     14'b00000010011101: fc_kernel = 8'h01;
     14'b00000010011110: fc_kernel = 8'h08;
     14'b00000010011111: fc_kernel = 8'h08;
     14'b00000010100000: fc_kernel = 8'h02;
     14'b00000010100001: fc_kernel = 8'h06;
     14'b00000010100010: fc_kernel = 8'h03;
     14'b00000010100011: fc_kernel = 8'h00;
     14'b00000010100100: fc_kernel = 8'h02;
     14'b00000010100101: fc_kernel = 8'h05;
     14'b00000010100110: fc_kernel = 8'hfd;
     14'b00000010100111: fc_kernel = 8'hc9;
     14'b00000010101000: fc_kernel = 8'h0d;
     14'b00000010101001: fc_kernel = 8'h03;
     14'b00000010101010: fc_kernel = 8'h07;
     14'b00000010101011: fc_kernel = 8'h01;
     14'b00000010101100: fc_kernel = 8'hf9;
     14'b00000010101101: fc_kernel = 8'hf4;
     14'b00000010101110: fc_kernel = 8'hfa;
     14'b00000010101111: fc_kernel = 8'hff;
     14'b00000010110000: fc_kernel = 8'hfd;
     14'b00000010110001: fc_kernel = 8'hfe;
     14'b00000010110010: fc_kernel = 8'hff;
     14'b00000010110011: fc_kernel = 8'h00;
     14'b00000010110100: fc_kernel = 8'h05;
     14'b00000010110101: fc_kernel = 8'h07;
     14'b00000010110110: fc_kernel = 8'h07;
     14'b00000010110111: fc_kernel = 8'h11;
     14'b00000010111000: fc_kernel = 8'h0d;
     14'b00000010111001: fc_kernel = 8'h08;
     14'b00000010111010: fc_kernel = 8'h02;
     14'b00000010111011: fc_kernel = 8'h00;
     14'b00000010111100: fc_kernel = 8'hfe;
     14'b00000010111101: fc_kernel = 8'h0a;
     14'b00000010111110: fc_kernel = 8'h08;
     14'b00000010111111: fc_kernel = 8'hd9;
     14'b00000011000000: fc_kernel = 8'h0c;
     14'b00000011000001: fc_kernel = 8'h03;
     14'b00000011000010: fc_kernel = 8'h05;
     14'b00000011000011: fc_kernel = 8'hfc;
     14'b00000011000100: fc_kernel = 8'hf8;
     14'b00000011000101: fc_kernel = 8'hf9;
     14'b00000011000110: fc_kernel = 8'hff;
     14'b00000011000111: fc_kernel = 8'hfd;
     14'b00000011001000: fc_kernel = 8'h00;
     14'b00000011001001: fc_kernel = 8'hf6;
     14'b00000011001010: fc_kernel = 8'h00;
     14'b00000011001011: fc_kernel = 8'h00;
     14'b00000011001100: fc_kernel = 8'hfc;
     14'b00000011001101: fc_kernel = 8'hfc;
     14'b00000011001110: fc_kernel = 8'hff;
     14'b00000011001111: fc_kernel = 8'h0a;
     14'b00000011010000: fc_kernel = 8'h05;
     14'b00000011010001: fc_kernel = 8'h09;
     14'b00000011010010: fc_kernel = 8'h00;
     14'b00000011010011: fc_kernel = 8'h00;
     14'b00000011010100: fc_kernel = 8'h00;
     14'b00000011010101: fc_kernel = 8'h05;
     14'b00000011010110: fc_kernel = 8'h00;
     14'b00000011010111: fc_kernel = 8'hda;
     14'b00000011011000: fc_kernel = 8'h0e;
     14'b00000011011001: fc_kernel = 8'hfc;
     14'b00000011011010: fc_kernel = 8'hfd;
     14'b00000011011011: fc_kernel = 8'hfa;
     14'b00000011011100: fc_kernel = 8'hf9;
     14'b00000011011101: fc_kernel = 8'hfb;
     14'b00000011011110: fc_kernel = 8'hfc;
     14'b00000011011111: fc_kernel = 8'hfa;
     14'b00000011100000: fc_kernel = 8'hfe;
     14'b00000011100001: fc_kernel = 8'hf7;
     14'b00000011100010: fc_kernel = 8'hfe;
     14'b00000011100011: fc_kernel = 8'hf8;
     14'b00000011100100: fc_kernel = 8'hf4;
     14'b00000011100101: fc_kernel = 8'he7;
     14'b00000011100110: fc_kernel = 8'hf2;
     14'b00000011100111: fc_kernel = 8'hff;
     14'b00000011101000: fc_kernel = 8'hfc;
     14'b00000011101001: fc_kernel = 8'h00;
     14'b00000011101010: fc_kernel = 8'h05;
     14'b00000011101011: fc_kernel = 8'h0b;
     14'b00000011101100: fc_kernel = 8'h09;
     14'b00000011101101: fc_kernel = 8'h09;
     14'b00000011101110: fc_kernel = 8'h00;
     14'b00000011101111: fc_kernel = 8'he3;
     14'b00000011110000: fc_kernel = 8'h05;
     14'b00000011110001: fc_kernel = 8'hfd;
     14'b00000011110010: fc_kernel = 8'hf8;
     14'b00000011110011: fc_kernel = 8'hff;
     14'b00000011110100: fc_kernel = 8'hff;
     14'b00000011110101: fc_kernel = 8'h00;
     14'b00000011110110: fc_kernel = 8'hfc;
     14'b00000011110111: fc_kernel = 8'hf6;
     14'b00000011111000: fc_kernel = 8'hfa;
     14'b00000011111001: fc_kernel = 8'hfe;
     14'b00000011111010: fc_kernel = 8'hfc;
     14'b00000011111011: fc_kernel = 8'hf8;
     14'b00000011111100: fc_kernel = 8'he3;
     14'b00000011111101: fc_kernel = 8'hdd;
     14'b00000011111110: fc_kernel = 8'hea;
     14'b00000011111111: fc_kernel = 8'hf9;
     14'b00000100000000: fc_kernel = 8'hfd;
     14'b00000100000001: fc_kernel = 8'hff;
     14'b00000100000010: fc_kernel = 8'hfe;
     14'b00000100000011: fc_kernel = 8'h0a;
     14'b00000100000100: fc_kernel = 8'h05;
     14'b00000100000101: fc_kernel = 8'h0e;
     14'b00000100000110: fc_kernel = 8'h09;
     14'b00000100000111: fc_kernel = 8'hf5;
     14'b00000100001000: fc_kernel = 8'h02;
     14'b00000100001001: fc_kernel = 8'hf6;
     14'b00000100001010: fc_kernel = 8'hf3;
     14'b00000100001011: fc_kernel = 8'h01;
     14'b00000100001100: fc_kernel = 8'h04;
     14'b00000100001101: fc_kernel = 8'h05;
     14'b00000100001110: fc_kernel = 8'h01;
     14'b00000100001111: fc_kernel = 8'hfc;
     14'b00000100010000: fc_kernel = 8'h00;
     14'b00000100010001: fc_kernel = 8'h03;
     14'b00000100010010: fc_kernel = 8'h00;
     14'b00000100010011: fc_kernel = 8'hf4;
     14'b00000100010100: fc_kernel = 8'hdf;
     14'b00000100010101: fc_kernel = 8'hdc;
     14'b00000100010110: fc_kernel = 8'he6;
     14'b00000100010111: fc_kernel = 8'hfa;
     14'b00000100011000: fc_kernel = 8'hfc;
     14'b00000100011001: fc_kernel = 8'hfb;
     14'b00000100011010: fc_kernel = 8'hfa;
     14'b00000100011011: fc_kernel = 8'hfe;
     14'b00000100011100: fc_kernel = 8'h02;
     14'b00000100011101: fc_kernel = 8'h0e;
     14'b00000100011110: fc_kernel = 8'h0c;
     14'b00000100011111: fc_kernel = 8'h08;
     14'b00000100100000: fc_kernel = 8'hf0;
     14'b00000100100001: fc_kernel = 8'hef;
     14'b00000100100010: fc_kernel = 8'hfc;
     14'b00000100100011: fc_kernel = 8'h03;
     14'b00000100100100: fc_kernel = 8'h09;
     14'b00000100100101: fc_kernel = 8'h06;
     14'b00000100100110: fc_kernel = 8'h09;
     14'b00000100100111: fc_kernel = 8'h06;
     14'b00000100101000: fc_kernel = 8'hfe;
     14'b00000100101001: fc_kernel = 8'h05;
     14'b00000100101010: fc_kernel = 8'h07;
     14'b00000100101011: fc_kernel = 8'hef;
     14'b00000100101100: fc_kernel = 8'hde;
     14'b00000100101101: fc_kernel = 8'hd4;
     14'b00000100101110: fc_kernel = 8'he2;
     14'b00000100101111: fc_kernel = 8'hf9;
     14'b00000100110000: fc_kernel = 8'h00;
     14'b00000100110001: fc_kernel = 8'hfb;
     14'b00000100110010: fc_kernel = 8'hfb;
     14'b00000100110011: fc_kernel = 8'hfe;
     14'b00000100110100: fc_kernel = 8'h03;
     14'b00000100110101: fc_kernel = 8'h0f;
     14'b00000100110110: fc_kernel = 8'h15;
     14'b00000100110111: fc_kernel = 8'h0e;
     14'b00000100111000: fc_kernel = 8'he9;
     14'b00000100111001: fc_kernel = 8'hf3;
     14'b00000100111010: fc_kernel = 8'h07;
     14'b00000100111011: fc_kernel = 8'h07;
     14'b00000100111100: fc_kernel = 8'h03;
     14'b00000100111101: fc_kernel = 8'h08;
     14'b00000100111110: fc_kernel = 8'h08;
     14'b00000100111111: fc_kernel = 8'h01;
     14'b00000101000000: fc_kernel = 8'h06;
     14'b00000101000001: fc_kernel = 8'h01;
     14'b00000101000010: fc_kernel = 8'hfb;
     14'b00000101000011: fc_kernel = 8'heb;
     14'b00000101000100: fc_kernel = 8'hda;
     14'b00000101000101: fc_kernel = 8'hd5;
     14'b00000101000110: fc_kernel = 8'he5;
     14'b00000101000111: fc_kernel = 8'hf4;
     14'b00000101001000: fc_kernel = 8'hf9;
     14'b00000101001001: fc_kernel = 8'hf7;
     14'b00000101001010: fc_kernel = 8'h02;
     14'b00000101001011: fc_kernel = 8'h06;
     14'b00000101001100: fc_kernel = 8'h08;
     14'b00000101001101: fc_kernel = 8'h0c;
     14'b00000101001110: fc_kernel = 8'h0c;
     14'b00000101001111: fc_kernel = 8'h05;
     14'b00000101010000: fc_kernel = 8'hf0;
     14'b00000101010001: fc_kernel = 8'hfd;
     14'b00000101010010: fc_kernel = 8'h0f;
     14'b00000101010011: fc_kernel = 8'h08;
     14'b00000101010100: fc_kernel = 8'h0c;
     14'b00000101010101: fc_kernel = 8'h0a;
     14'b00000101010110: fc_kernel = 8'h0d;
     14'b00000101010111: fc_kernel = 8'h09;
     14'b00000101011000: fc_kernel = 8'h05;
     14'b00000101011001: fc_kernel = 8'h05;
     14'b00000101011010: fc_kernel = 8'hf8;
     14'b00000101011011: fc_kernel = 8'hdc;
     14'b00000101011100: fc_kernel = 8'hd5;
     14'b00000101011101: fc_kernel = 8'hde;
     14'b00000101011110: fc_kernel = 8'hec;
     14'b00000101011111: fc_kernel = 8'hfb;
     14'b00000101100000: fc_kernel = 8'hfd;
     14'b00000101100001: fc_kernel = 8'h03;
     14'b00000101100010: fc_kernel = 8'h08;
     14'b00000101100011: fc_kernel = 8'h03;
     14'b00000101100100: fc_kernel = 8'h00;
     14'b00000101100101: fc_kernel = 8'h0a;
     14'b00000101100110: fc_kernel = 8'h03;
     14'b00000101100111: fc_kernel = 8'hfa;
     14'b00000101101000: fc_kernel = 8'he2;
     14'b00000101101001: fc_kernel = 8'hfa;
     14'b00000101101010: fc_kernel = 8'h0a;
     14'b00000101101011: fc_kernel = 8'h05;
     14'b00000101101100: fc_kernel = 8'h08;
     14'b00000101101101: fc_kernel = 8'h01;
     14'b00000101101110: fc_kernel = 8'h0c;
     14'b00000101101111: fc_kernel = 8'h0e;
     14'b00000101110000: fc_kernel = 8'h10;
     14'b00000101110001: fc_kernel = 8'h07;
     14'b00000101110010: fc_kernel = 8'hef;
     14'b00000101110011: fc_kernel = 8'hd8;
     14'b00000101110100: fc_kernel = 8'hda;
     14'b00000101110101: fc_kernel = 8'heb;
     14'b00000101110110: fc_kernel = 8'hfd;
     14'b00000101110111: fc_kernel = 8'h03;
     14'b00000101111000: fc_kernel = 8'h02;
     14'b00000101111001: fc_kernel = 8'hff;
     14'b00000101111010: fc_kernel = 8'h06;
     14'b00000101111011: fc_kernel = 8'h03;
     14'b00000101111100: fc_kernel = 8'h02;
     14'b00000101111101: fc_kernel = 8'h04;
     14'b00000101111110: fc_kernel = 8'hff;
     14'b00000101111111: fc_kernel = 8'hf3;
     14'b00000110000000: fc_kernel = 8'he7;
     14'b00000110000001: fc_kernel = 8'hf9;
     14'b00000110000010: fc_kernel = 8'hff;
     14'b00000110000011: fc_kernel = 8'h01;
     14'b00000110000100: fc_kernel = 8'h03;
     14'b00000110000101: fc_kernel = 8'h03;
     14'b00000110000110: fc_kernel = 8'h08;
     14'b00000110000111: fc_kernel = 8'h0e;
     14'b00000110001000: fc_kernel = 8'h14;
     14'b00000110001001: fc_kernel = 8'h09;
     14'b00000110001010: fc_kernel = 8'hf3;
     14'b00000110001011: fc_kernel = 8'hde;
     14'b00000110001100: fc_kernel = 8'he3;
     14'b00000110001101: fc_kernel = 8'hf4;
     14'b00000110001110: fc_kernel = 8'h00;
     14'b00000110001111: fc_kernel = 8'h01;
     14'b00000110010000: fc_kernel = 8'h05;
     14'b00000110010001: fc_kernel = 8'h03;
     14'b00000110010010: fc_kernel = 8'h00;
     14'b00000110010011: fc_kernel = 8'h06;
     14'b00000110010100: fc_kernel = 8'h04;
     14'b00000110010101: fc_kernel = 8'h08;
     14'b00000110010110: fc_kernel = 8'hfd;
     14'b00000110010111: fc_kernel = 8'hf4;
     14'b00000110011000: fc_kernel = 8'hee;
     14'b00000110011001: fc_kernel = 8'hf4;
     14'b00000110011010: fc_kernel = 8'h00;
     14'b00000110011011: fc_kernel = 8'h04;
     14'b00000110011100: fc_kernel = 8'h00;
     14'b00000110011101: fc_kernel = 8'h09;
     14'b00000110011110: fc_kernel = 8'h0b;
     14'b00000110011111: fc_kernel = 8'h0f;
     14'b00000110100000: fc_kernel = 8'h0e;
     14'b00000110100001: fc_kernel = 8'h0f;
     14'b00000110100010: fc_kernel = 8'h00;
     14'b00000110100011: fc_kernel = 8'hed;
     14'b00000110100100: fc_kernel = 8'hef;
     14'b00000110100101: fc_kernel = 8'hf6;
     14'b00000110100110: fc_kernel = 8'hfe;
     14'b00000110100111: fc_kernel = 8'h03;
     14'b00000110101000: fc_kernel = 8'h01;
     14'b00000110101001: fc_kernel = 8'h01;
     14'b00000110101010: fc_kernel = 8'h00;
     14'b00000110101011: fc_kernel = 8'h05;
     14'b00000110101100: fc_kernel = 8'h09;
     14'b00000110101101: fc_kernel = 8'h00;
     14'b00000110101110: fc_kernel = 8'hfa;
     14'b00000110101111: fc_kernel = 8'hfb;
     14'b00000110110000: fc_kernel = 8'hed;
     14'b00000110110001: fc_kernel = 8'hfc;
     14'b00000110110010: fc_kernel = 8'h01;
     14'b00000110110011: fc_kernel = 8'h08;
     14'b00000110110100: fc_kernel = 8'h04;
     14'b00000110110101: fc_kernel = 8'h09;
     14'b00000110110110: fc_kernel = 8'h03;
     14'b00000110110111: fc_kernel = 8'h07;
     14'b00000110111000: fc_kernel = 8'h0d;
     14'b00000110111001: fc_kernel = 8'h0c;
     14'b00000110111010: fc_kernel = 8'h08;
     14'b00000110111011: fc_kernel = 8'hfb;
     14'b00000110111100: fc_kernel = 8'hf9;
     14'b00000110111101: fc_kernel = 8'hfd;
     14'b00000110111110: fc_kernel = 8'hff;
     14'b00000110111111: fc_kernel = 8'h00;
     14'b00000111000000: fc_kernel = 8'hfe;
     14'b00000111000001: fc_kernel = 8'hfa;
     14'b00000111000010: fc_kernel = 8'hfe;
     14'b00000111000011: fc_kernel = 8'h05;
     14'b00000111000100: fc_kernel = 8'h05;
     14'b00000111000101: fc_kernel = 8'h00;
     14'b00000111000110: fc_kernel = 8'hf5;
     14'b00000111000111: fc_kernel = 8'hf2;
     14'b00000111001000: fc_kernel = 8'hf8;
     14'b00000111001001: fc_kernel = 8'hfd;
     14'b00000111001010: fc_kernel = 8'hfd;
     14'b00000111001011: fc_kernel = 8'h08;
     14'b00000111001100: fc_kernel = 8'h03;
     14'b00000111001101: fc_kernel = 8'h00;
     14'b00000111001110: fc_kernel = 8'h04;
     14'b00000111001111: fc_kernel = 8'h03;
     14'b00000111010000: fc_kernel = 8'h06;
     14'b00000111010001: fc_kernel = 8'h10;
     14'b00000111010010: fc_kernel = 8'h08;
     14'b00000111010011: fc_kernel = 8'h04;
     14'b00000111010100: fc_kernel = 8'h01;
     14'b00000111010101: fc_kernel = 8'hfd;
     14'b00000111010110: fc_kernel = 8'h01;
     14'b00000111010111: fc_kernel = 8'hff;
     14'b00000111011000: fc_kernel = 8'hfc;
     14'b00000111011001: fc_kernel = 8'hfc;
     14'b00000111011010: fc_kernel = 8'hfc;
     14'b00000111011011: fc_kernel = 8'h01;
     14'b00000111011100: fc_kernel = 8'h05;
     14'b00000111011101: fc_kernel = 8'hf9;
     14'b00000111011110: fc_kernel = 8'hf4;
     14'b00000111011111: fc_kernel = 8'hee;
     14'b00000111100000: fc_kernel = 8'hfa;
     14'b00000111100001: fc_kernel = 8'hf4;
     14'b00000111100010: fc_kernel = 8'hf6;
     14'b00000111100011: fc_kernel = 8'h00;
     14'b00000111100100: fc_kernel = 8'h06;
     14'b00000111100101: fc_kernel = 8'h08;
     14'b00000111100110: fc_kernel = 8'h04;
     14'b00000111100111: fc_kernel = 8'h0a;
     14'b00000111101000: fc_kernel = 8'h09;
     14'b00000111101001: fc_kernel = 8'h0e;
     14'b00000111101010: fc_kernel = 8'h09;
     14'b00000111101011: fc_kernel = 8'h09;
     14'b00000111101100: fc_kernel = 8'h00;
     14'b00000111101101: fc_kernel = 8'h00;
     14'b00000111101110: fc_kernel = 8'h04;
     14'b00000111101111: fc_kernel = 8'hfa;
     14'b00000111110000: fc_kernel = 8'hfd;
     14'b00000111110001: fc_kernel = 8'hfb;
     14'b00000111110010: fc_kernel = 8'hfc;
     14'b00000111110011: fc_kernel = 8'h04;
     14'b00000111110100: fc_kernel = 8'h00;
     14'b00000111110101: fc_kernel = 8'h02;
     14'b00000111110110: fc_kernel = 8'hf8;
     14'b00000111110111: fc_kernel = 8'hee;
     14'b00000111111000: fc_kernel = 8'hf8;
     14'b00000111111001: fc_kernel = 8'heb;
     14'b00000111111010: fc_kernel = 8'hf1;
     14'b00000111111011: fc_kernel = 8'hf9;
     14'b00000111111100: fc_kernel = 8'hfe;
     14'b00000111111101: fc_kernel = 8'h01;
     14'b00000111111110: fc_kernel = 8'h07;
     14'b00000111111111: fc_kernel = 8'h10;
     14'b00001000000000: fc_kernel = 8'h0f;
     14'b00001000000001: fc_kernel = 8'h0e;
     14'b00001000000010: fc_kernel = 8'h10;
     14'b00001000000011: fc_kernel = 8'h12;
     14'b00001000000100: fc_kernel = 8'h10;
     14'b00001000000101: fc_kernel = 8'h09;
     14'b00001000000110: fc_kernel = 8'h05;
     14'b00001000000111: fc_kernel = 8'h06;
     14'b00001000001000: fc_kernel = 8'h00;
     14'b00001000001001: fc_kernel = 8'hfb;
     14'b00001000001010: fc_kernel = 8'hf7;
     14'b00001000001011: fc_kernel = 8'hfd;
     14'b00001000001100: fc_kernel = 8'h03;
     14'b00001000001101: fc_kernel = 8'h00;
     14'b00001000001110: fc_kernel = 8'hf3;
     14'b00001000001111: fc_kernel = 8'hf0;
     14'b00001000010000: fc_kernel = 8'hef;
     14'b00001000010001: fc_kernel = 8'he6;
     14'b00001000010010: fc_kernel = 8'hef;
     14'b00001000010011: fc_kernel = 8'hf9;
     14'b00001000010100: fc_kernel = 8'hff;
     14'b00001000010101: fc_kernel = 8'hff;
     14'b00001000010110: fc_kernel = 8'h00;
     14'b00001000010111: fc_kernel = 8'h02;
     14'b00001000011000: fc_kernel = 8'h06;
     14'b00001000011001: fc_kernel = 8'h04;
     14'b00001000011010: fc_kernel = 8'h0c;
     14'b00001000011011: fc_kernel = 8'h08;
     14'b00001000011100: fc_kernel = 8'h05;
     14'b00001000011101: fc_kernel = 8'hfe;
     14'b00001000011110: fc_kernel = 8'h00;
     14'b00001000011111: fc_kernel = 8'hf8;
     14'b00001000100000: fc_kernel = 8'hf3;
     14'b00001000100001: fc_kernel = 8'he7;
     14'b00001000100010: fc_kernel = 8'heb;
     14'b00001000100011: fc_kernel = 8'hee;
     14'b00001000100100: fc_kernel = 8'hf4;
     14'b00001000100101: fc_kernel = 8'heb;
     14'b00001000100110: fc_kernel = 8'he8;
     14'b00001000100111: fc_kernel = 8'heb;
     14'b00001000101000: fc_kernel = 8'he4;
     14'b00001000101001: fc_kernel = 8'hd9;
     14'b00001000101010: fc_kernel = 8'hed;
     14'b00001000101011: fc_kernel = 8'hf3;
     14'b00001000101100: fc_kernel = 8'hf1;
     14'b00001000101101: fc_kernel = 8'hea;
     14'b00001000101110: fc_kernel = 8'hed;
     14'b00001000101111: fc_kernel = 8'heb;
     14'b00001000110000: fc_kernel = 8'heb;
     14'b00001000110001: fc_kernel = 8'he7;
     14'b00001000110010: fc_kernel = 8'he9;
     14'b00001000110011: fc_kernel = 8'hec;
     14'b00001000110100: fc_kernel = 8'he7;
     14'b00001000110101: fc_kernel = 8'hdf;
     14'b00001000110110: fc_kernel = 8'he4;
     14'b00001000110111: fc_kernel = 8'he2;
     14'b00001000111000: fc_kernel = 8'hd9;
     14'b00001000111001: fc_kernel = 8'hcf;
     14'b00001000111010: fc_kernel = 8'hcd;
     14'b00001000111011: fc_kernel = 8'hd0;
     14'b00001000111100: fc_kernel = 8'hd9;
     14'b00001000111101: fc_kernel = 8'hd9;
     14'b00001000111110: fc_kernel = 8'hde;
     14'b00001000111111: fc_kernel = 8'he6;
     14'b00010000000000: fc_kernel = 8'h0d;
     14'b00010000000001: fc_kernel = 8'h0b;
     14'b00010000000010: fc_kernel = 8'he6;
     14'b00010000000011: fc_kernel = 8'hfb;
     14'b00010000000100: fc_kernel = 8'h11;
     14'b00010000000101: fc_kernel = 8'hf4;
     14'b00010000000110: fc_kernel = 8'hf3;
     14'b00010000000111: fc_kernel = 8'hf3;
     14'b00010000001000: fc_kernel = 8'hfb;
     14'b00010000001001: fc_kernel = 8'h0c;
     14'b00010000001010: fc_kernel = 8'h16;
     14'b00010000001011: fc_kernel = 8'h0b;
     14'b00010000001100: fc_kernel = 8'h0b;
     14'b00010000001101: fc_kernel = 8'h1c;
     14'b00010000001110: fc_kernel = 8'h1f;
     14'b00010000001111: fc_kernel = 8'h0d;
     14'b00010000010000: fc_kernel = 8'h02;
     14'b00010000010001: fc_kernel = 8'h00;
     14'b00010000010010: fc_kernel = 8'h01;
     14'b00010000010011: fc_kernel = 8'hf5;
     14'b00010000010100: fc_kernel = 8'hf6;
     14'b00010000010101: fc_kernel = 8'hfc;
     14'b00010000010110: fc_kernel = 8'hff;
     14'b00010000010111: fc_kernel = 8'hfe;
     14'b00010000011000: fc_kernel = 8'h14;
     14'b00010000011001: fc_kernel = 8'h11;
     14'b00010000011010: fc_kernel = 8'h07;
     14'b00010000011011: fc_kernel = 8'hf7;
     14'b00010000011100: fc_kernel = 8'hf5;
     14'b00010000011101: fc_kernel = 8'hfe;
     14'b00010000011110: fc_kernel = 8'hf3;
     14'b00010000011111: fc_kernel = 8'hf0;
     14'b00010000100000: fc_kernel = 8'he9;
     14'b00010000100001: fc_kernel = 8'hf0;
     14'b00010000100010: fc_kernel = 8'hfb;
     14'b00010000100011: fc_kernel = 8'hfb;
     14'b00010000100100: fc_kernel = 8'hf3;
     14'b00010000100101: fc_kernel = 8'h01;
     14'b00010000100110: fc_kernel = 8'h08;
     14'b00010000100111: fc_kernel = 8'hfa;
     14'b00010000101000: fc_kernel = 8'hef;
     14'b00010000101001: fc_kernel = 8'hf0;
     14'b00010000101010: fc_kernel = 8'hf4;
     14'b00010000101011: fc_kernel = 8'hec;
     14'b00010000101100: fc_kernel = 8'he8;
     14'b00010000101101: fc_kernel = 8'he4;
     14'b00010000101110: fc_kernel = 8'he5;
     14'b00010000101111: fc_kernel = 8'he7;
     14'b00010000110000: fc_kernel = 8'h17;
     14'b00010000110001: fc_kernel = 8'hfd;
     14'b00010000110010: fc_kernel = 8'h0b;
     14'b00010000110011: fc_kernel = 8'h09;
     14'b00010000110100: fc_kernel = 8'hff;
     14'b00010000110101: fc_kernel = 8'h03;
     14'b00010000110110: fc_kernel = 8'hfc;
     14'b00010000110111: fc_kernel = 8'hfe;
     14'b00010000111000: fc_kernel = 8'hed;
     14'b00010000111001: fc_kernel = 8'heb;
     14'b00010000111010: fc_kernel = 8'hf3;
     14'b00010000111011: fc_kernel = 8'hfb;
     14'b00010000111100: fc_kernel = 8'hf7;
     14'b00010000111101: fc_kernel = 8'hf6;
     14'b00010000111110: fc_kernel = 8'hfb;
     14'b00010000111111: fc_kernel = 8'hf0;
     14'b00010001000000: fc_kernel = 8'hef;
     14'b00010001000001: fc_kernel = 8'hf1;
     14'b00010001000010: fc_kernel = 8'hf7;
     14'b00010001000011: fc_kernel = 8'hf3;
     14'b00010001000100: fc_kernel = 8'he8;
     14'b00010001000101: fc_kernel = 8'he3;
     14'b00010001000110: fc_kernel = 8'hdd;
     14'b00010001000111: fc_kernel = 8'hd1;
     14'b00010001001000: fc_kernel = 8'h19;
     14'b00010001001001: fc_kernel = 8'h04;
     14'b00010001001010: fc_kernel = 8'h13;
     14'b00010001001011: fc_kernel = 8'h14;
     14'b00010001001100: fc_kernel = 8'h09;
     14'b00010001001101: fc_kernel = 8'h04;
     14'b00010001001110: fc_kernel = 8'hf3;
     14'b00010001001111: fc_kernel = 8'hf1;
     14'b00010001010000: fc_kernel = 8'hf2;
     14'b00010001010001: fc_kernel = 8'hf0;
     14'b00010001010010: fc_kernel = 8'hf1;
     14'b00010001010011: fc_kernel = 8'hf7;
     14'b00010001010100: fc_kernel = 8'hf8;
     14'b00010001010101: fc_kernel = 8'hf9;
     14'b00010001010110: fc_kernel = 8'hf4;
     14'b00010001010111: fc_kernel = 8'heb;
     14'b00010001011000: fc_kernel = 8'hf2;
     14'b00010001011001: fc_kernel = 8'hf6;
     14'b00010001011010: fc_kernel = 8'hf5;
     14'b00010001011011: fc_kernel = 8'hfc;
     14'b00010001011100: fc_kernel = 8'hfa;
     14'b00010001011101: fc_kernel = 8'h00;
     14'b00010001011110: fc_kernel = 8'hf4;
     14'b00010001011111: fc_kernel = 8'hd9;
     14'b00010001100000: fc_kernel = 8'hfe;
     14'b00010001100001: fc_kernel = 8'h09;
     14'b00010001100010: fc_kernel = 8'h09;
     14'b00010001100011: fc_kernel = 8'h07;
     14'b00010001100100: fc_kernel = 8'h01;
     14'b00010001100101: fc_kernel = 8'hf6;
     14'b00010001100110: fc_kernel = 8'hf0;
     14'b00010001100111: fc_kernel = 8'hf4;
     14'b00010001101000: fc_kernel = 8'hf7;
     14'b00010001101001: fc_kernel = 8'hf1;
     14'b00010001101010: fc_kernel = 8'hf0;
     14'b00010001101011: fc_kernel = 8'hf5;
     14'b00010001101100: fc_kernel = 8'hf9;
     14'b00010001101101: fc_kernel = 8'hf6;
     14'b00010001101110: fc_kernel = 8'hed;
     14'b00010001101111: fc_kernel = 8'hf1;
     14'b00010001110000: fc_kernel = 8'hf2;
     14'b00010001110001: fc_kernel = 8'hfd;
     14'b00010001110010: fc_kernel = 8'hfc;
     14'b00010001110011: fc_kernel = 8'h01;
     14'b00010001110100: fc_kernel = 8'h02;
     14'b00010001110101: fc_kernel = 8'h02;
     14'b00010001110110: fc_kernel = 8'hf9;
     14'b00010001110111: fc_kernel = 8'hde;
     14'b00010001111000: fc_kernel = 8'heb;
     14'b00010001111001: fc_kernel = 8'hfe;
     14'b00010001111010: fc_kernel = 8'h06;
     14'b00010001111011: fc_kernel = 8'hfb;
     14'b00010001111100: fc_kernel = 8'hf0;
     14'b00010001111101: fc_kernel = 8'hef;
     14'b00010001111110: fc_kernel = 8'hed;
     14'b00010001111111: fc_kernel = 8'hef;
     14'b00010010000000: fc_kernel = 8'hf5;
     14'b00010010000001: fc_kernel = 8'hf3;
     14'b00010010000010: fc_kernel = 8'hf9;
     14'b00010010000011: fc_kernel = 8'hf8;
     14'b00010010000100: fc_kernel = 8'hf3;
     14'b00010010000101: fc_kernel = 8'hf1;
     14'b00010010000110: fc_kernel = 8'heb;
     14'b00010010000111: fc_kernel = 8'hec;
     14'b00010010001000: fc_kernel = 8'hf4;
     14'b00010010001001: fc_kernel = 8'hfb;
     14'b00010010001010: fc_kernel = 8'hfe;
     14'b00010010001011: fc_kernel = 8'hfd;
     14'b00010010001100: fc_kernel = 8'hfb;
     14'b00010010001101: fc_kernel = 8'hf5;
     14'b00010010001110: fc_kernel = 8'hea;
     14'b00010010001111: fc_kernel = 8'hcb;
     14'b00010010010000: fc_kernel = 8'he6;
     14'b00010010010001: fc_kernel = 8'hee;
     14'b00010010010010: fc_kernel = 8'hf2;
     14'b00010010010011: fc_kernel = 8'hed;
     14'b00010010010100: fc_kernel = 8'hf3;
     14'b00010010010101: fc_kernel = 8'hf0;
     14'b00010010010110: fc_kernel = 8'hef;
     14'b00010010010111: fc_kernel = 8'hf1;
     14'b00010010011000: fc_kernel = 8'hf5;
     14'b00010010011001: fc_kernel = 8'hf2;
     14'b00010010011010: fc_kernel = 8'hf4;
     14'b00010010011011: fc_kernel = 8'hfa;
     14'b00010010011100: fc_kernel = 8'hfd;
     14'b00010010011101: fc_kernel = 8'hf1;
     14'b00010010011110: fc_kernel = 8'hf1;
     14'b00010010011111: fc_kernel = 8'hf6;
     14'b00010010100000: fc_kernel = 8'hf8;
     14'b00010010100001: fc_kernel = 8'hfa;
     14'b00010010100010: fc_kernel = 8'hfc;
     14'b00010010100011: fc_kernel = 8'hfc;
     14'b00010010100100: fc_kernel = 8'hf3;
     14'b00010010100101: fc_kernel = 8'he9;
     14'b00010010100110: fc_kernel = 8'hdf;
     14'b00010010100111: fc_kernel = 8'hc1;
     14'b00010010101000: fc_kernel = 8'hda;
     14'b00010010101001: fc_kernel = 8'hea;
     14'b00010010101010: fc_kernel = 8'he5;
     14'b00010010101011: fc_kernel = 8'he3;
     14'b00010010101100: fc_kernel = 8'hf4;
     14'b00010010101101: fc_kernel = 8'hfd;
     14'b00010010101110: fc_kernel = 8'hfa;
     14'b00010010101111: fc_kernel = 8'hee;
     14'b00010010110000: fc_kernel = 8'hfb;
     14'b00010010110001: fc_kernel = 8'hfd;
     14'b00010010110010: fc_kernel = 8'hff;
     14'b00010010110011: fc_kernel = 8'h02;
     14'b00010010110100: fc_kernel = 8'h03;
     14'b00010010110101: fc_kernel = 8'h07;
     14'b00010010110110: fc_kernel = 8'hfe;
     14'b00010010110111: fc_kernel = 8'hfe;
     14'b00010010111000: fc_kernel = 8'hff;
     14'b00010010111001: fc_kernel = 8'hf6;
     14'b00010010111010: fc_kernel = 8'hf2;
     14'b00010010111011: fc_kernel = 8'hf0;
     14'b00010010111100: fc_kernel = 8'hf4;
     14'b00010010111101: fc_kernel = 8'he5;
     14'b00010010111110: fc_kernel = 8'hd9;
     14'b00010010111111: fc_kernel = 8'hce;
     14'b00010011000000: fc_kernel = 8'he5;
     14'b00010011000001: fc_kernel = 8'hec;
     14'b00010011000010: fc_kernel = 8'he7;
     14'b00010011000011: fc_kernel = 8'hd7;
     14'b00010011000100: fc_kernel = 8'hdf;
     14'b00010011000101: fc_kernel = 8'hf5;
     14'b00010011000110: fc_kernel = 8'hf2;
     14'b00010011000111: fc_kernel = 8'hf3;
     14'b00010011001000: fc_kernel = 8'hfc;
     14'b00010011001001: fc_kernel = 8'hfd;
     14'b00010011001010: fc_kernel = 8'h00;
     14'b00010011001011: fc_kernel = 8'h00;
     14'b00010011001100: fc_kernel = 8'h10;
     14'b00010011001101: fc_kernel = 8'h13;
     14'b00010011001110: fc_kernel = 8'h0b;
     14'b00010011001111: fc_kernel = 8'hfe;
     14'b00010011010000: fc_kernel = 8'hfd;
     14'b00010011010001: fc_kernel = 8'hef;
     14'b00010011010010: fc_kernel = 8'hf4;
     14'b00010011010011: fc_kernel = 8'hf4;
     14'b00010011010100: fc_kernel = 8'hf6;
     14'b00010011010101: fc_kernel = 8'he2;
     14'b00010011010110: fc_kernel = 8'hd6;
     14'b00010011010111: fc_kernel = 8'hd3;
     14'b00010011011000: fc_kernel = 8'heb;
     14'b00010011011001: fc_kernel = 8'hf1;
     14'b00010011011010: fc_kernel = 8'he9;
     14'b00010011011011: fc_kernel = 8'he3;
     14'b00010011011100: fc_kernel = 8'he3;
     14'b00010011011101: fc_kernel = 8'hf0;
     14'b00010011011110: fc_kernel = 8'hed;
     14'b00010011011111: fc_kernel = 8'hf1;
     14'b00010011100000: fc_kernel = 8'hf9;
     14'b00010011100001: fc_kernel = 8'hfc;
     14'b00010011100010: fc_kernel = 8'hfb;
     14'b00010011100011: fc_kernel = 8'h09;
     14'b00010011100100: fc_kernel = 8'h1d;
     14'b00010011100101: fc_kernel = 8'h1b;
     14'b00010011100110: fc_kernel = 8'h0c;
     14'b00010011100111: fc_kernel = 8'hfd;
     14'b00010011101000: fc_kernel = 8'hf4;
     14'b00010011101001: fc_kernel = 8'hf8;
     14'b00010011101010: fc_kernel = 8'hf4;
     14'b00010011101011: fc_kernel = 8'hf9;
     14'b00010011101100: fc_kernel = 8'hf8;
     14'b00010011101101: fc_kernel = 8'hed;
     14'b00010011101110: fc_kernel = 8'he3;
     14'b00010011101111: fc_kernel = 8'hdb;
     14'b00010011110000: fc_kernel = 8'hef;
     14'b00010011110001: fc_kernel = 8'hfa;
     14'b00010011110010: fc_kernel = 8'hef;
     14'b00010011110011: fc_kernel = 8'hed;
     14'b00010011110100: fc_kernel = 8'hf5;
     14'b00010011110101: fc_kernel = 8'hf5;
     14'b00010011110110: fc_kernel = 8'hfa;
     14'b00010011110111: fc_kernel = 8'hf4;
     14'b00010011111000: fc_kernel = 8'hf3;
     14'b00010011111001: fc_kernel = 8'hf5;
     14'b00010011111010: fc_kernel = 8'hfb;
     14'b00010011111011: fc_kernel = 8'h0f;
     14'b00010011111100: fc_kernel = 8'h1f;
     14'b00010011111101: fc_kernel = 8'h17;
     14'b00010011111110: fc_kernel = 8'h0a;
     14'b00010011111111: fc_kernel = 8'h01;
     14'b00010100000000: fc_kernel = 8'hf6;
     14'b00010100000001: fc_kernel = 8'hf6;
     14'b00010100000010: fc_kernel = 8'hf6;
     14'b00010100000011: fc_kernel = 8'h00;
     14'b00010100000100: fc_kernel = 8'hff;
     14'b00010100000101: fc_kernel = 8'hfe;
     14'b00010100000110: fc_kernel = 8'hf0;
     14'b00010100000111: fc_kernel = 8'he5;
     14'b00010100001000: fc_kernel = 8'hfa;
     14'b00010100001001: fc_kernel = 8'h08;
     14'b00010100001010: fc_kernel = 8'h00;
     14'b00010100001011: fc_kernel = 8'hfb;
     14'b00010100001100: fc_kernel = 8'hf8;
     14'b00010100001101: fc_kernel = 8'hfd;
     14'b00010100001110: fc_kernel = 8'hfd;
     14'b00010100001111: fc_kernel = 8'hfd;
     14'b00010100010000: fc_kernel = 8'hec;
     14'b00010100010001: fc_kernel = 8'he5;
     14'b00010100010010: fc_kernel = 8'hfa;
     14'b00010100010011: fc_kernel = 8'h0f;
     14'b00010100010100: fc_kernel = 8'h21;
     14'b00010100010101: fc_kernel = 8'h14;
     14'b00010100010110: fc_kernel = 8'h10;
     14'b00010100010111: fc_kernel = 8'h00;
     14'b00010100011000: fc_kernel = 8'hf6;
     14'b00010100011001: fc_kernel = 8'hf4;
     14'b00010100011010: fc_kernel = 8'hf6;
     14'b00010100011011: fc_kernel = 8'hff;
     14'b00010100011100: fc_kernel = 8'h03;
     14'b00010100011101: fc_kernel = 8'hf3;
     14'b00010100011110: fc_kernel = 8'hf2;
     14'b00010100011111: fc_kernel = 8'he3;
     14'b00010100100000: fc_kernel = 8'h0d;
     14'b00010100100001: fc_kernel = 8'h18;
     14'b00010100100010: fc_kernel = 8'h0c;
     14'b00010100100011: fc_kernel = 8'h00;
     14'b00010100100100: fc_kernel = 8'hf5;
     14'b00010100100101: fc_kernel = 8'hfb;
     14'b00010100100110: fc_kernel = 8'h00;
     14'b00010100100111: fc_kernel = 8'hf5;
     14'b00010100101000: fc_kernel = 8'hdd;
     14'b00010100101001: fc_kernel = 8'he7;
     14'b00010100101010: fc_kernel = 8'h03;
     14'b00010100101011: fc_kernel = 8'h19;
     14'b00010100101100: fc_kernel = 8'h1d;
     14'b00010100101101: fc_kernel = 8'h18;
     14'b00010100101110: fc_kernel = 8'h09;
     14'b00010100101111: fc_kernel = 8'hfe;
     14'b00010100110000: fc_kernel = 8'hea;
     14'b00010100110001: fc_kernel = 8'he8;
     14'b00010100110010: fc_kernel = 8'hf2;
     14'b00010100110011: fc_kernel = 8'hf9;
     14'b00010100110100: fc_kernel = 8'hfb;
     14'b00010100110101: fc_kernel = 8'hfb;
     14'b00010100110110: fc_kernel = 8'hf6;
     14'b00010100110111: fc_kernel = 8'hf3;
     14'b00010100111000: fc_kernel = 8'h19;
     14'b00010100111001: fc_kernel = 8'h15;
     14'b00010100111010: fc_kernel = 8'hff;
     14'b00010100111011: fc_kernel = 8'hef;
     14'b00010100111100: fc_kernel = 8'hee;
     14'b00010100111101: fc_kernel = 8'hfa;
     14'b00010100111110: fc_kernel = 8'h06;
     14'b00010100111111: fc_kernel = 8'hf1;
     14'b00010101000000: fc_kernel = 8'he9;
     14'b00010101000001: fc_kernel = 8'heb;
     14'b00010101000010: fc_kernel = 8'h04;
     14'b00010101000011: fc_kernel = 8'h1e;
     14'b00010101000100: fc_kernel = 8'h19;
     14'b00010101000101: fc_kernel = 8'h15;
     14'b00010101000110: fc_kernel = 8'h06;
     14'b00010101000111: fc_kernel = 8'hf3;
     14'b00010101001000: fc_kernel = 8'he2;
     14'b00010101001001: fc_kernel = 8'hd9;
     14'b00010101001010: fc_kernel = 8'he1;
     14'b00010101001011: fc_kernel = 8'he8;
     14'b00010101001100: fc_kernel = 8'hf2;
     14'b00010101001101: fc_kernel = 8'hed;
     14'b00010101001110: fc_kernel = 8'hf1;
     14'b00010101001111: fc_kernel = 8'hf1;
     14'b00010101010000: fc_kernel = 8'h14;
     14'b00010101010001: fc_kernel = 8'h03;
     14'b00010101010010: fc_kernel = 8'hf3;
     14'b00010101010011: fc_kernel = 8'hed;
     14'b00010101010100: fc_kernel = 8'hec;
     14'b00010101010101: fc_kernel = 8'hfb;
     14'b00010101010110: fc_kernel = 8'hfd;
     14'b00010101010111: fc_kernel = 8'hf6;
     14'b00010101011000: fc_kernel = 8'hec;
     14'b00010101011001: fc_kernel = 8'hf2;
     14'b00010101011010: fc_kernel = 8'h0b;
     14'b00010101011011: fc_kernel = 8'h1e;
     14'b00010101011100: fc_kernel = 8'h15;
     14'b00010101011101: fc_kernel = 8'h16;
     14'b00010101011110: fc_kernel = 8'hf6;
     14'b00010101011111: fc_kernel = 8'he4;
     14'b00010101100000: fc_kernel = 8'hd8;
     14'b00010101100001: fc_kernel = 8'hd9;
     14'b00010101100010: fc_kernel = 8'he5;
     14'b00010101100011: fc_kernel = 8'hf6;
     14'b00010101100100: fc_kernel = 8'hf4;
     14'b00010101100101: fc_kernel = 8'hed;
     14'b00010101100110: fc_kernel = 8'hec;
     14'b00010101100111: fc_kernel = 8'he8;
     14'b00010101101000: fc_kernel = 8'hef;
     14'b00010101101001: fc_kernel = 8'hd3;
     14'b00010101101010: fc_kernel = 8'hea;
     14'b00010101101011: fc_kernel = 8'hde;
     14'b00010101101100: fc_kernel = 8'hde;
     14'b00010101101101: fc_kernel = 8'hf3;
     14'b00010101101110: fc_kernel = 8'hfb;
     14'b00010101101111: fc_kernel = 8'hfb;
     14'b00010101110000: fc_kernel = 8'hef;
     14'b00010101110001: fc_kernel = 8'hf5;
     14'b00010101110010: fc_kernel = 8'h08;
     14'b00010101110011: fc_kernel = 8'h1c;
     14'b00010101110100: fc_kernel = 8'h18;
     14'b00010101110101: fc_kernel = 8'h0d;
     14'b00010101110110: fc_kernel = 8'he6;
     14'b00010101110111: fc_kernel = 8'hda;
     14'b00010101111000: fc_kernel = 8'hda;
     14'b00010101111001: fc_kernel = 8'hf0;
     14'b00010101111010: fc_kernel = 8'h00;
     14'b00010101111011: fc_kernel = 8'h01;
     14'b00010101111100: fc_kernel = 8'hff;
     14'b00010101111101: fc_kernel = 8'hfb;
     14'b00010101111110: fc_kernel = 8'hf4;
     14'b00010101111111: fc_kernel = 8'heb;
     14'b00010110000000: fc_kernel = 8'hfa;
     14'b00010110000001: fc_kernel = 8'hdc;
     14'b00010110000010: fc_kernel = 8'he2;
     14'b00010110000011: fc_kernel = 8'hc9;
     14'b00010110000100: fc_kernel = 8'hdb;
     14'b00010110000101: fc_kernel = 8'hec;
     14'b00010110000110: fc_kernel = 8'hf4;
     14'b00010110000111: fc_kernel = 8'hfa;
     14'b00010110001000: fc_kernel = 8'hf3;
     14'b00010110001001: fc_kernel = 8'hf1;
     14'b00010110001010: fc_kernel = 8'h0b;
     14'b00010110001011: fc_kernel = 8'h13;
     14'b00010110001100: fc_kernel = 8'h12;
     14'b00010110001101: fc_kernel = 8'h05;
     14'b00010110001110: fc_kernel = 8'he2;
     14'b00010110001111: fc_kernel = 8'he1;
     14'b00010110010000: fc_kernel = 8'hf2;
     14'b00010110010001: fc_kernel = 8'hfd;
     14'b00010110010010: fc_kernel = 8'h01;
     14'b00010110010011: fc_kernel = 8'h04;
     14'b00010110010100: fc_kernel = 8'hfb;
     14'b00010110010101: fc_kernel = 8'hfd;
     14'b00010110010110: fc_kernel = 8'hfc;
     14'b00010110010111: fc_kernel = 8'h03;
     14'b00010110011000: fc_kernel = 8'h0b;
     14'b00010110011001: fc_kernel = 8'h0c;
     14'b00010110011010: fc_kernel = 8'hc4;
     14'b00010110011011: fc_kernel = 8'hcc;
     14'b00010110011100: fc_kernel = 8'he6;
     14'b00010110011101: fc_kernel = 8'hfc;
     14'b00010110011110: fc_kernel = 8'h00;
     14'b00010110011111: fc_kernel = 8'h01;
     14'b00010110100000: fc_kernel = 8'hfa;
     14'b00010110100001: fc_kernel = 8'hfa;
     14'b00010110100010: fc_kernel = 8'h08;
     14'b00010110100011: fc_kernel = 8'h11;
     14'b00010110100100: fc_kernel = 8'h06;
     14'b00010110100101: fc_kernel = 8'hff;
     14'b00010110100110: fc_kernel = 8'hf3;
     14'b00010110100111: fc_kernel = 8'hf9;
     14'b00010110101000: fc_kernel = 8'h07;
     14'b00010110101001: fc_kernel = 8'h0f;
     14'b00010110101010: fc_kernel = 8'h0a;
     14'b00010110101011: fc_kernel = 8'h05;
     14'b00010110101100: fc_kernel = 8'h01;
     14'b00010110101101: fc_kernel = 8'h00;
     14'b00010110101110: fc_kernel = 8'h04;
     14'b00010110101111: fc_kernel = 8'h0d;
     14'b00010110110000: fc_kernel = 8'h0b;
     14'b00010110110001: fc_kernel = 8'h14;
     14'b00010110110010: fc_kernel = 8'hd1;
     14'b00010110110011: fc_kernel = 8'hda;
     14'b00010110110100: fc_kernel = 8'hf2;
     14'b00010110110101: fc_kernel = 8'h00;
     14'b00010110110110: fc_kernel = 8'h06;
     14'b00010110110111: fc_kernel = 8'h06;
     14'b00010110111000: fc_kernel = 8'h05;
     14'b00010110111001: fc_kernel = 8'h02;
     14'b00010110111010: fc_kernel = 8'h0a;
     14'b00010110111011: fc_kernel = 8'h08;
     14'b00010110111100: fc_kernel = 8'h04;
     14'b00010110111101: fc_kernel = 8'h03;
     14'b00010110111110: fc_kernel = 8'h00;
     14'b00010110111111: fc_kernel = 8'h0a;
     14'b00010111000000: fc_kernel = 8'h0f;
     14'b00010111000001: fc_kernel = 8'h0b;
     14'b00010111000010: fc_kernel = 8'h06;
     14'b00010111000011: fc_kernel = 8'h02;
     14'b00010111000100: fc_kernel = 8'h00;
     14'b00010111000101: fc_kernel = 8'hfd;
     14'b00010111000110: fc_kernel = 8'h05;
     14'b00010111000111: fc_kernel = 8'h0e;
     14'b00010111001000: fc_kernel = 8'h00;
     14'b00010111001001: fc_kernel = 8'h0b;
     14'b00010111001010: fc_kernel = 8'h0c;
     14'b00010111001011: fc_kernel = 8'h0b;
     14'b00010111001100: fc_kernel = 8'h06;
     14'b00010111001101: fc_kernel = 8'h06;
     14'b00010111001110: fc_kernel = 8'h05;
     14'b00010111001111: fc_kernel = 8'h06;
     14'b00010111010000: fc_kernel = 8'h05;
     14'b00010111010001: fc_kernel = 8'h00;
     14'b00010111010010: fc_kernel = 8'hf7;
     14'b00010111010011: fc_kernel = 8'hff;
     14'b00010111010100: fc_kernel = 8'h00;
     14'b00010111010101: fc_kernel = 8'hff;
     14'b00010111010110: fc_kernel = 8'h00;
     14'b00010111010111: fc_kernel = 8'h07;
     14'b00010111011000: fc_kernel = 8'h11;
     14'b00010111011001: fc_kernel = 8'h11;
     14'b00010111011010: fc_kernel = 8'h0e;
     14'b00010111011011: fc_kernel = 8'h06;
     14'b00010111011100: fc_kernel = 8'hff;
     14'b00010111011101: fc_kernel = 8'hfa;
     14'b00010111011110: fc_kernel = 8'h05;
     14'b00010111011111: fc_kernel = 8'h14;
     14'b00010111100000: fc_kernel = 8'hf1;
     14'b00010111100001: fc_kernel = 8'h00;
     14'b00010111100010: fc_kernel = 8'h0e;
     14'b00010111100011: fc_kernel = 8'h1e;
     14'b00010111100100: fc_kernel = 8'h12;
     14'b00010111100101: fc_kernel = 8'h07;
     14'b00010111100110: fc_kernel = 8'h06;
     14'b00010111100111: fc_kernel = 8'h06;
     14'b00010111101000: fc_kernel = 8'h00;
     14'b00010111101001: fc_kernel = 8'h01;
     14'b00010111101010: fc_kernel = 8'hf9;
     14'b00010111101011: fc_kernel = 8'hf8;
     14'b00010111101100: fc_kernel = 8'hfe;
     14'b00010111101101: fc_kernel = 8'h06;
     14'b00010111101110: fc_kernel = 8'h05;
     14'b00010111101111: fc_kernel = 8'h0a;
     14'b00010111110000: fc_kernel = 8'h07;
     14'b00010111110001: fc_kernel = 8'h0d;
     14'b00010111110010: fc_kernel = 8'h09;
     14'b00010111110011: fc_kernel = 8'h01;
     14'b00010111110100: fc_kernel = 8'hfc;
     14'b00010111110101: fc_kernel = 8'hf3;
     14'b00010111110110: fc_kernel = 8'h00;
     14'b00010111110111: fc_kernel = 8'h13;
     14'b00010111111000: fc_kernel = 8'hf6;
     14'b00010111111001: fc_kernel = 8'hf5;
     14'b00010111111010: fc_kernel = 8'h0a;
     14'b00010111111011: fc_kernel = 8'h19;
     14'b00010111111100: fc_kernel = 8'h12;
     14'b00010111111101: fc_kernel = 8'h05;
     14'b00010111111110: fc_kernel = 8'h00;
     14'b00010111111111: fc_kernel = 8'h07;
     14'b00011000000000: fc_kernel = 8'h01;
     14'b00011000000001: fc_kernel = 8'h00;
     14'b00011000000010: fc_kernel = 8'hfd;
     14'b00011000000011: fc_kernel = 8'hff;
     14'b00011000000100: fc_kernel = 8'hfc;
     14'b00011000000101: fc_kernel = 8'h01;
     14'b00011000000110: fc_kernel = 8'h0a;
     14'b00011000000111: fc_kernel = 8'h07;
     14'b00011000001000: fc_kernel = 8'h0b;
     14'b00011000001001: fc_kernel = 8'h0c;
     14'b00011000001010: fc_kernel = 8'h04;
     14'b00011000001011: fc_kernel = 8'hfb;
     14'b00011000001100: fc_kernel = 8'hee;
     14'b00011000001101: fc_kernel = 8'hee;
     14'b00011000001110: fc_kernel = 8'hf4;
     14'b00011000001111: fc_kernel = 8'h0c;
     14'b00011000010000: fc_kernel = 8'hf7;
     14'b00011000010001: fc_kernel = 8'hf7;
     14'b00011000010010: fc_kernel = 8'hfc;
     14'b00011000010011: fc_kernel = 8'h04;
     14'b00011000010100: fc_kernel = 8'h03;
     14'b00011000010101: fc_kernel = 8'hfb;
     14'b00011000010110: fc_kernel = 8'hfb;
     14'b00011000010111: fc_kernel = 8'hfb;
     14'b00011000011000: fc_kernel = 8'hf3;
     14'b00011000011001: fc_kernel = 8'hf4;
     14'b00011000011010: fc_kernel = 8'hf6;
     14'b00011000011011: fc_kernel = 8'hf9;
     14'b00011000011100: fc_kernel = 8'hf5;
     14'b00011000011101: fc_kernel = 8'hf3;
     14'b00011000011110: fc_kernel = 8'hfa;
     14'b00011000011111: fc_kernel = 8'h00;
     14'b00011000100000: fc_kernel = 8'h08;
     14'b00011000100001: fc_kernel = 8'h06;
     14'b00011000100010: fc_kernel = 8'h05;
     14'b00011000100011: fc_kernel = 8'hf5;
     14'b00011000100100: fc_kernel = 8'hef;
     14'b00011000100101: fc_kernel = 8'he9;
     14'b00011000100110: fc_kernel = 8'hee;
     14'b00011000100111: fc_kernel = 8'h0a;
     14'b00011000101000: fc_kernel = 8'he7;
     14'b00011000101001: fc_kernel = 8'heb;
     14'b00011000101010: fc_kernel = 8'hef;
     14'b00011000101011: fc_kernel = 8'hf4;
     14'b00011000101100: fc_kernel = 8'hed;
     14'b00011000101101: fc_kernel = 8'hef;
     14'b00011000101110: fc_kernel = 8'hf8;
     14'b00011000101111: fc_kernel = 8'hea;
     14'b00011000110000: fc_kernel = 8'he2;
     14'b00011000110001: fc_kernel = 8'he3;
     14'b00011000110010: fc_kernel = 8'he8;
     14'b00011000110011: fc_kernel = 8'he9;
     14'b00011000110100: fc_kernel = 8'he9;
     14'b00011000110101: fc_kernel = 8'hd9;
     14'b00011000110110: fc_kernel = 8'hda;
     14'b00011000110111: fc_kernel = 8'hd9;
     14'b00011000111000: fc_kernel = 8'hf1;
     14'b00011000111001: fc_kernel = 8'hfe;
     14'b00011000111010: fc_kernel = 8'hfa;
     14'b00011000111011: fc_kernel = 8'hf2;
     14'b00011000111100: fc_kernel = 8'hf4;
     14'b00011000111101: fc_kernel = 8'he5;
     14'b00011000111110: fc_kernel = 8'hef;
     14'b00011000111111: fc_kernel = 8'h04;
     14'b00100000000000: fc_kernel = 8'he9;
     14'b00100000000001: fc_kernel = 8'h04;
     14'b00100000000010: fc_kernel = 8'h04;
     14'b00100000000011: fc_kernel = 8'he8;
     14'b00100000000100: fc_kernel = 8'hf7;
     14'b00100000000101: fc_kernel = 8'h09;
     14'b00100000000110: fc_kernel = 8'h10;
     14'b00100000000111: fc_kernel = 8'h11;
     14'b00100000001000: fc_kernel = 8'h17;
     14'b00100000001001: fc_kernel = 8'h11;
     14'b00100000001010: fc_kernel = 8'h16;
     14'b00100000001011: fc_kernel = 8'h09;
     14'b00100000001100: fc_kernel = 8'h0e;
     14'b00100000001101: fc_kernel = 8'h0c;
     14'b00100000001110: fc_kernel = 8'h09;
     14'b00100000001111: fc_kernel = 8'h01;
     14'b00100000010000: fc_kernel = 8'hf4;
     14'b00100000010001: fc_kernel = 8'hec;
     14'b00100000010010: fc_kernel = 8'hee;
     14'b00100000010011: fc_kernel = 8'hf4;
     14'b00100000010100: fc_kernel = 8'he5;
     14'b00100000010101: fc_kernel = 8'hfe;
     14'b00100000010110: fc_kernel = 8'h0a;
     14'b00100000010111: fc_kernel = 8'h0d;
     14'b00100000011000: fc_kernel = 8'h00;
     14'b00100000011001: fc_kernel = 8'hf7;
     14'b00100000011010: fc_kernel = 8'hf1;
     14'b00100000011011: fc_kernel = 8'hef;
     14'b00100000011100: fc_kernel = 8'h00;
     14'b00100000011101: fc_kernel = 8'h03;
     14'b00100000011110: fc_kernel = 8'h1b;
     14'b00100000011111: fc_kernel = 8'h16;
     14'b00100000100000: fc_kernel = 8'h19;
     14'b00100000100001: fc_kernel = 8'h1b;
     14'b00100000100010: fc_kernel = 8'h16;
     14'b00100000100011: fc_kernel = 8'h12;
     14'b00100000100100: fc_kernel = 8'h11;
     14'b00100000100101: fc_kernel = 8'h0d;
     14'b00100000100110: fc_kernel = 8'h0a;
     14'b00100000100111: fc_kernel = 8'h02;
     14'b00100000101000: fc_kernel = 8'hfb;
     14'b00100000101001: fc_kernel = 8'hf9;
     14'b00100000101010: fc_kernel = 8'hf6;
     14'b00100000101011: fc_kernel = 8'hf4;
     14'b00100000101100: fc_kernel = 8'hef;
     14'b00100000101101: fc_kernel = 8'heb;
     14'b00100000101110: fc_kernel = 8'h04;
     14'b00100000101111: fc_kernel = 8'h09;
     14'b00100000110000: fc_kernel = 8'h08;
     14'b00100000110001: fc_kernel = 8'hea;
     14'b00100000110010: fc_kernel = 8'hfa;
     14'b00100000110011: fc_kernel = 8'h06;
     14'b00100000110100: fc_kernel = 8'h0c;
     14'b00100000110101: fc_kernel = 8'h0c;
     14'b00100000110110: fc_kernel = 8'h12;
     14'b00100000110111: fc_kernel = 8'h14;
     14'b00100000111000: fc_kernel = 8'h15;
     14'b00100000111001: fc_kernel = 8'h0f;
     14'b00100000111010: fc_kernel = 8'h0a;
     14'b00100000111011: fc_kernel = 8'h0b;
     14'b00100000111100: fc_kernel = 8'h08;
     14'b00100000111101: fc_kernel = 8'h06;
     14'b00100000111110: fc_kernel = 8'h06;
     14'b00100000111111: fc_kernel = 8'h04;
     14'b00100001000000: fc_kernel = 8'hff;
     14'b00100001000001: fc_kernel = 8'hfe;
     14'b00100001000010: fc_kernel = 8'h00;
     14'b00100001000011: fc_kernel = 8'hf4;
     14'b00100001000100: fc_kernel = 8'he9;
     14'b00100001000101: fc_kernel = 8'he4;
     14'b00100001000110: fc_kernel = 8'hf5;
     14'b00100001000111: fc_kernel = 8'hff;
     14'b00100001001000: fc_kernel = 8'h00;
     14'b00100001001001: fc_kernel = 8'h00;
     14'b00100001001010: fc_kernel = 8'h00;
     14'b00100001001011: fc_kernel = 8'hfd;
     14'b00100001001100: fc_kernel = 8'h08;
     14'b00100001001101: fc_kernel = 8'h03;
     14'b00100001001110: fc_kernel = 8'h02;
     14'b00100001001111: fc_kernel = 8'h05;
     14'b00100001010000: fc_kernel = 8'h03;
     14'b00100001010001: fc_kernel = 8'h07;
     14'b00100001010010: fc_kernel = 8'h05;
     14'b00100001010011: fc_kernel = 8'h00;
     14'b00100001010100: fc_kernel = 8'h08;
     14'b00100001010101: fc_kernel = 8'h08;
     14'b00100001010110: fc_kernel = 8'h07;
     14'b00100001010111: fc_kernel = 8'h0d;
     14'b00100001011000: fc_kernel = 8'h01;
     14'b00100001011001: fc_kernel = 8'h00;
     14'b00100001011010: fc_kernel = 8'h02;
     14'b00100001011011: fc_kernel = 8'h00;
     14'b00100001011100: fc_kernel = 8'hfb;
     14'b00100001011101: fc_kernel = 8'hee;
     14'b00100001011110: fc_kernel = 8'he6;
     14'b00100001011111: fc_kernel = 8'hef;
     14'b00100001100000: fc_kernel = 8'h03;
     14'b00100001100001: fc_kernel = 8'h08;
     14'b00100001100010: fc_kernel = 8'h04;
     14'b00100001100011: fc_kernel = 8'h06;
     14'b00100001100100: fc_kernel = 8'h02;
     14'b00100001100101: fc_kernel = 8'h07;
     14'b00100001100110: fc_kernel = 8'h0a;
     14'b00100001100111: fc_kernel = 8'h01;
     14'b00100001101000: fc_kernel = 8'h02;
     14'b00100001101001: fc_kernel = 8'h05;
     14'b00100001101010: fc_kernel = 8'h04;
     14'b00100001101011: fc_kernel = 8'h04;
     14'b00100001101100: fc_kernel = 8'h04;
     14'b00100001101101: fc_kernel = 8'h03;
     14'b00100001101110: fc_kernel = 8'h07;
     14'b00100001101111: fc_kernel = 8'h02;
     14'b00100001110000: fc_kernel = 8'h00;
     14'b00100001110001: fc_kernel = 8'h00;
     14'b00100001110010: fc_kernel = 8'hfa;
     14'b00100001110011: fc_kernel = 8'h01;
     14'b00100001110100: fc_kernel = 8'hfa;
     14'b00100001110101: fc_kernel = 8'hec;
     14'b00100001110110: fc_kernel = 8'hda;
     14'b00100001110111: fc_kernel = 8'hdf;
     14'b00100001111000: fc_kernel = 8'hff;
     14'b00100001111001: fc_kernel = 8'h0f;
     14'b00100001111010: fc_kernel = 8'h0b;
     14'b00100001111011: fc_kernel = 8'h03;
     14'b00100001111100: fc_kernel = 8'h04;
     14'b00100001111101: fc_kernel = 8'h00;
     14'b00100001111110: fc_kernel = 8'h04;
     14'b00100001111111: fc_kernel = 8'h04;
     14'b00100010000000: fc_kernel = 8'h04;
     14'b00100010000001: fc_kernel = 8'h02;
     14'b00100010000010: fc_kernel = 8'h00;
     14'b00100010000011: fc_kernel = 8'h03;
     14'b00100010000100: fc_kernel = 8'h04;
     14'b00100010000101: fc_kernel = 8'h05;
     14'b00100010000110: fc_kernel = 8'hfe;
     14'b00100010000111: fc_kernel = 8'hff;
     14'b00100010001000: fc_kernel = 8'hfd;
     14'b00100010001001: fc_kernel = 8'hfb;
     14'b00100010001010: fc_kernel = 8'hfb;
     14'b00100010001011: fc_kernel = 8'hff;
     14'b00100010001100: fc_kernel = 8'hfd;
     14'b00100010001101: fc_kernel = 8'hee;
     14'b00100010001110: fc_kernel = 8'hd2;
     14'b00100010001111: fc_kernel = 8'hdb;
     14'b00100010010000: fc_kernel = 8'hf6;
     14'b00100010010001: fc_kernel = 8'h0d;
     14'b00100010010010: fc_kernel = 8'h0d;
     14'b00100010010011: fc_kernel = 8'h05;
     14'b00100010010100: fc_kernel = 8'hfa;
     14'b00100010010101: fc_kernel = 8'h00;
     14'b00100010010110: fc_kernel = 8'hfc;
     14'b00100010010111: fc_kernel = 8'h02;
     14'b00100010011000: fc_kernel = 8'hfe;
     14'b00100010011001: fc_kernel = 8'h02;
     14'b00100010011010: fc_kernel = 8'h01;
     14'b00100010011011: fc_kernel = 8'h00;
     14'b00100010011100: fc_kernel = 8'h04;
     14'b00100010011101: fc_kernel = 8'h07;
     14'b00100010011110: fc_kernel = 8'hfd;
     14'b00100010011111: fc_kernel = 8'hff;
     14'b00100010100000: fc_kernel = 8'hff;
     14'b00100010100001: fc_kernel = 8'h01;
     14'b00100010100010: fc_kernel = 8'h00;
     14'b00100010100011: fc_kernel = 8'h00;
     14'b00100010100100: fc_kernel = 8'h00;
     14'b00100010100101: fc_kernel = 8'hfc;
     14'b00100010100110: fc_kernel = 8'he1;
     14'b00100010100111: fc_kernel = 8'hcb;
     14'b00100010101000: fc_kernel = 8'h01;
     14'b00100010101001: fc_kernel = 8'h07;
     14'b00100010101010: fc_kernel = 8'h04;
     14'b00100010101011: fc_kernel = 8'h07;
     14'b00100010101100: fc_kernel = 8'h00;
     14'b00100010101101: fc_kernel = 8'hfa;
     14'b00100010101110: fc_kernel = 8'hfe;
     14'b00100010101111: fc_kernel = 8'h05;
     14'b00100010110000: fc_kernel = 8'h05;
     14'b00100010110001: fc_kernel = 8'h04;
     14'b00100010110010: fc_kernel = 8'h00;
     14'b00100010110011: fc_kernel = 8'hff;
     14'b00100010110100: fc_kernel = 8'h09;
     14'b00100010110101: fc_kernel = 8'h06;
     14'b00100010110110: fc_kernel = 8'h09;
     14'b00100010110111: fc_kernel = 8'h02;
     14'b00100010111000: fc_kernel = 8'h03;
     14'b00100010111001: fc_kernel = 8'h01;
     14'b00100010111010: fc_kernel = 8'hff;
     14'b00100010111011: fc_kernel = 8'hfc;
     14'b00100010111100: fc_kernel = 8'hff;
     14'b00100010111101: fc_kernel = 8'hf8;
     14'b00100010111110: fc_kernel = 8'he6;
     14'b00100010111111: fc_kernel = 8'hbe;
     14'b00100011000000: fc_kernel = 8'hff;
     14'b00100011000001: fc_kernel = 8'h03;
     14'b00100011000010: fc_kernel = 8'h06;
     14'b00100011000011: fc_kernel = 8'h0a;
     14'b00100011000100: fc_kernel = 8'h06;
     14'b00100011000101: fc_kernel = 8'h00;
     14'b00100011000110: fc_kernel = 8'hfe;
     14'b00100011000111: fc_kernel = 8'h00;
     14'b00100011001000: fc_kernel = 8'h03;
     14'b00100011001001: fc_kernel = 8'hfe;
     14'b00100011001010: fc_kernel = 8'hff;
     14'b00100011001011: fc_kernel = 8'hfe;
     14'b00100011001100: fc_kernel = 8'h00;
     14'b00100011001101: fc_kernel = 8'h00;
     14'b00100011001110: fc_kernel = 8'h00;
     14'b00100011001111: fc_kernel = 8'h03;
     14'b00100011010000: fc_kernel = 8'h01;
     14'b00100011010001: fc_kernel = 8'h00;
     14'b00100011010010: fc_kernel = 8'h01;
     14'b00100011010011: fc_kernel = 8'hf8;
     14'b00100011010100: fc_kernel = 8'hfe;
     14'b00100011010101: fc_kernel = 8'hfa;
     14'b00100011010110: fc_kernel = 8'he5;
     14'b00100011010111: fc_kernel = 8'hd4;
     14'b00100011011000: fc_kernel = 8'hfa;
     14'b00100011011001: fc_kernel = 8'h01;
     14'b00100011011010: fc_kernel = 8'h09;
     14'b00100011011011: fc_kernel = 8'h0e;
     14'b00100011011100: fc_kernel = 8'h06;
     14'b00100011011101: fc_kernel = 8'hfe;
     14'b00100011011110: fc_kernel = 8'hfb;
     14'b00100011011111: fc_kernel = 8'hf5;
     14'b00100011100000: fc_kernel = 8'hec;
     14'b00100011100001: fc_kernel = 8'heb;
     14'b00100011100010: fc_kernel = 8'hea;
     14'b00100011100011: fc_kernel = 8'hde;
     14'b00100011100100: fc_kernel = 8'he2;
     14'b00100011100101: fc_kernel = 8'hec;
     14'b00100011100110: fc_kernel = 8'hf2;
     14'b00100011100111: fc_kernel = 8'hfa;
     14'b00100011101000: fc_kernel = 8'h00;
     14'b00100011101001: fc_kernel = 8'h02;
     14'b00100011101010: fc_kernel = 8'h02;
     14'b00100011101011: fc_kernel = 8'h00;
     14'b00100011101100: fc_kernel = 8'hfe;
     14'b00100011101101: fc_kernel = 8'hf8;
     14'b00100011101110: fc_kernel = 8'hf4;
     14'b00100011101111: fc_kernel = 8'hf9;
     14'b00100011110000: fc_kernel = 8'hfb;
     14'b00100011110001: fc_kernel = 8'hfa;
     14'b00100011110010: fc_kernel = 8'hfd;
     14'b00100011110011: fc_kernel = 8'hf9;
     14'b00100011110100: fc_kernel = 8'he8;
     14'b00100011110101: fc_kernel = 8'he5;
     14'b00100011110110: fc_kernel = 8'he4;
     14'b00100011110111: fc_kernel = 8'hed;
     14'b00100011111000: fc_kernel = 8'he5;
     14'b00100011111001: fc_kernel = 8'he5;
     14'b00100011111010: fc_kernel = 8'hdf;
     14'b00100011111011: fc_kernel = 8'hdf;
     14'b00100011111100: fc_kernel = 8'hde;
     14'b00100011111101: fc_kernel = 8'he8;
     14'b00100011111110: fc_kernel = 8'hf3;
     14'b00100011111111: fc_kernel = 8'hf1;
     14'b00100100000000: fc_kernel = 8'hf7;
     14'b00100100000001: fc_kernel = 8'hf9;
     14'b00100100000010: fc_kernel = 8'hfd;
     14'b00100100000011: fc_kernel = 8'hfa;
     14'b00100100000100: fc_kernel = 8'hf9;
     14'b00100100000101: fc_kernel = 8'hf0;
     14'b00100100000110: fc_kernel = 8'h02;
     14'b00100100000111: fc_kernel = 8'h23;
     14'b00100100001000: fc_kernel = 8'hfb;
     14'b00100100001001: fc_kernel = 8'hec;
     14'b00100100001010: fc_kernel = 8'hd9;
     14'b00100100001011: fc_kernel = 8'hd7;
     14'b00100100001100: fc_kernel = 8'hd1;
     14'b00100100001101: fc_kernel = 8'hd9;
     14'b00100100001110: fc_kernel = 8'he5;
     14'b00100100001111: fc_kernel = 8'heb;
     14'b00100100010000: fc_kernel = 8'hf0;
     14'b00100100010001: fc_kernel = 8'hf7;
     14'b00100100010010: fc_kernel = 8'hfa;
     14'b00100100010011: fc_kernel = 8'hfd;
     14'b00100100010100: fc_kernel = 8'hf8;
     14'b00100100010101: fc_kernel = 8'hf1;
     14'b00100100010110: fc_kernel = 8'hf2;
     14'b00100100010111: fc_kernel = 8'hf9;
     14'b00100100011000: fc_kernel = 8'hfd;
     14'b00100100011001: fc_kernel = 8'h00;
     14'b00100100011010: fc_kernel = 8'hff;
     14'b00100100011011: fc_kernel = 8'hfe;
     14'b00100100011100: fc_kernel = 8'hf6;
     14'b00100100011101: fc_kernel = 8'hfa;
     14'b00100100011110: fc_kernel = 8'h0c;
     14'b00100100011111: fc_kernel = 8'h40;
     14'b00100100100000: fc_kernel = 8'hfa;
     14'b00100100100001: fc_kernel = 8'he7;
     14'b00100100100010: fc_kernel = 8'hd1;
     14'b00100100100011: fc_kernel = 8'hd2;
     14'b00100100100100: fc_kernel = 8'hd9;
     14'b00100100100101: fc_kernel = 8'hed;
     14'b00100100100110: fc_kernel = 8'hf5;
     14'b00100100100111: fc_kernel = 8'hf7;
     14'b00100100101000: fc_kernel = 8'hf8;
     14'b00100100101001: fc_kernel = 8'hfe;
     14'b00100100101010: fc_kernel = 8'hfd;
     14'b00100100101011: fc_kernel = 8'hfd;
     14'b00100100101100: fc_kernel = 8'hff;
     14'b00100100101101: fc_kernel = 8'hf6;
     14'b00100100101110: fc_kernel = 8'hf7;
     14'b00100100101111: fc_kernel = 8'hf9;
     14'b00100100110000: fc_kernel = 8'hf9;
     14'b00100100110001: fc_kernel = 8'h00;
     14'b00100100110010: fc_kernel = 8'hf9;
     14'b00100100110011: fc_kernel = 8'hf9;
     14'b00100100110100: fc_kernel = 8'hfb;
     14'b00100100110101: fc_kernel = 8'h01;
     14'b00100100110110: fc_kernel = 8'h14;
     14'b00100100110111: fc_kernel = 8'h35;
     14'b00100100111000: fc_kernel = 8'hfb;
     14'b00100100111001: fc_kernel = 8'hf7;
     14'b00100100111010: fc_kernel = 8'hed;
     14'b00100100111011: fc_kernel = 8'hf8;
     14'b00100100111100: fc_kernel = 8'hf3;
     14'b00100100111101: fc_kernel = 8'hfc;
     14'b00100100111110: fc_kernel = 8'hf8;
     14'b00100100111111: fc_kernel = 8'hfa;
     14'b00100101000000: fc_kernel = 8'hfd;
     14'b00100101000001: fc_kernel = 8'hf4;
     14'b00100101000010: fc_kernel = 8'hf9;
     14'b00100101000011: fc_kernel = 8'h05;
     14'b00100101000100: fc_kernel = 8'hfd;
     14'b00100101000101: fc_kernel = 8'hfd;
     14'b00100101000110: fc_kernel = 8'h00;
     14'b00100101000111: fc_kernel = 8'hf9;
     14'b00100101001000: fc_kernel = 8'hfd;
     14'b00100101001001: fc_kernel = 8'hfb;
     14'b00100101001010: fc_kernel = 8'h00;
     14'b00100101001011: fc_kernel = 8'hf7;
     14'b00100101001100: fc_kernel = 8'hf9;
     14'b00100101001101: fc_kernel = 8'hfd;
     14'b00100101001110: fc_kernel = 8'h16;
     14'b00100101001111: fc_kernel = 8'h37;
     14'b00100101010000: fc_kernel = 8'h07;
     14'b00100101010001: fc_kernel = 8'h0c;
     14'b00100101010010: fc_kernel = 8'h08;
     14'b00100101010011: fc_kernel = 8'h09;
     14'b00100101010100: fc_kernel = 8'h07;
     14'b00100101010101: fc_kernel = 8'hf9;
     14'b00100101010110: fc_kernel = 8'hfe;
     14'b00100101010111: fc_kernel = 8'h00;
     14'b00100101011000: fc_kernel = 8'h01;
     14'b00100101011001: fc_kernel = 8'h05;
     14'b00100101011010: fc_kernel = 8'h04;
     14'b00100101011011: fc_kernel = 8'h09;
     14'b00100101011100: fc_kernel = 8'h02;
     14'b00100101011101: fc_kernel = 8'hfe;
     14'b00100101011110: fc_kernel = 8'h03;
     14'b00100101011111: fc_kernel = 8'hff;
     14'b00100101100000: fc_kernel = 8'h02;
     14'b00100101100001: fc_kernel = 8'hff;
     14'b00100101100010: fc_kernel = 8'h00;
     14'b00100101100011: fc_kernel = 8'h04;
     14'b00100101100100: fc_kernel = 8'h00;
     14'b00100101100101: fc_kernel = 8'hfe;
     14'b00100101100110: fc_kernel = 8'h0f;
     14'b00100101100111: fc_kernel = 8'h38;
     14'b00100101101000: fc_kernel = 8'h0e;
     14'b00100101101001: fc_kernel = 8'h0f;
     14'b00100101101010: fc_kernel = 8'h12;
     14'b00100101101011: fc_kernel = 8'h0f;
     14'b00100101101100: fc_kernel = 8'h06;
     14'b00100101101101: fc_kernel = 8'h01;
     14'b00100101101110: fc_kernel = 8'hfd;
     14'b00100101101111: fc_kernel = 8'hfe;
     14'b00100101110000: fc_kernel = 8'h02;
     14'b00100101110001: fc_kernel = 8'h05;
     14'b00100101110010: fc_kernel = 8'h09;
     14'b00100101110011: fc_kernel = 8'h0b;
     14'b00100101110100: fc_kernel = 8'h02;
     14'b00100101110101: fc_kernel = 8'hff;
     14'b00100101110110: fc_kernel = 8'h00;
     14'b00100101110111: fc_kernel = 8'hfe;
     14'b00100101111000: fc_kernel = 8'h02;
     14'b00100101111001: fc_kernel = 8'hfc;
     14'b00100101111010: fc_kernel = 8'h01;
     14'b00100101111011: fc_kernel = 8'h01;
     14'b00100101111100: fc_kernel = 8'h02;
     14'b00100101111101: fc_kernel = 8'h02;
     14'b00100101111110: fc_kernel = 8'h15;
     14'b00100101111111: fc_kernel = 8'h39;
     14'b00100110000000: fc_kernel = 8'h0a;
     14'b00100110000001: fc_kernel = 8'h09;
     14'b00100110000010: fc_kernel = 8'h12;
     14'b00100110000011: fc_kernel = 8'h0b;
     14'b00100110000100: fc_kernel = 8'h00;
     14'b00100110000101: fc_kernel = 8'h00;
     14'b00100110000110: fc_kernel = 8'hff;
     14'b00100110000111: fc_kernel = 8'h03;
     14'b00100110001000: fc_kernel = 8'h03;
     14'b00100110001001: fc_kernel = 8'h09;
     14'b00100110001010: fc_kernel = 8'h0e;
     14'b00100110001011: fc_kernel = 8'h0e;
     14'b00100110001100: fc_kernel = 8'h05;
     14'b00100110001101: fc_kernel = 8'h01;
     14'b00100110001110: fc_kernel = 8'h07;
     14'b00100110001111: fc_kernel = 8'h0b;
     14'b00100110010000: fc_kernel = 8'h06;
     14'b00100110010001: fc_kernel = 8'h00;
     14'b00100110010010: fc_kernel = 8'hfe;
     14'b00100110010011: fc_kernel = 8'h02;
     14'b00100110010100: fc_kernel = 8'h0c;
     14'b00100110010101: fc_kernel = 8'h04;
     14'b00100110010110: fc_kernel = 8'h14;
     14'b00100110010111: fc_kernel = 8'h38;
     14'b00100110011000: fc_kernel = 8'hf8;
     14'b00100110011001: fc_kernel = 8'h02;
     14'b00100110011010: fc_kernel = 8'h0b;
     14'b00100110011011: fc_kernel = 8'h05;
     14'b00100110011100: fc_kernel = 8'h02;
     14'b00100110011101: fc_kernel = 8'h05;
     14'b00100110011110: fc_kernel = 8'h08;
     14'b00100110011111: fc_kernel = 8'h02;
     14'b00100110100000: fc_kernel = 8'h0a;
     14'b00100110100001: fc_kernel = 8'h06;
     14'b00100110100010: fc_kernel = 8'h0a;
     14'b00100110100011: fc_kernel = 8'h0c;
     14'b00100110100100: fc_kernel = 8'h02;
     14'b00100110100101: fc_kernel = 8'h05;
     14'b00100110100110: fc_kernel = 8'h03;
     14'b00100110100111: fc_kernel = 8'h07;
     14'b00100110101000: fc_kernel = 8'h01;
     14'b00100110101001: fc_kernel = 8'h00;
     14'b00100110101010: fc_kernel = 8'h00;
     14'b00100110101011: fc_kernel = 8'h06;
     14'b00100110101100: fc_kernel = 8'h06;
     14'b00100110101101: fc_kernel = 8'h03;
     14'b00100110101110: fc_kernel = 8'h15;
     14'b00100110101111: fc_kernel = 8'h27;
     14'b00100110110000: fc_kernel = 8'hfd;
     14'b00100110110001: fc_kernel = 8'h04;
     14'b00100110110010: fc_kernel = 8'h02;
     14'b00100110110011: fc_kernel = 8'h01;
     14'b00100110110100: fc_kernel = 8'h08;
     14'b00100110110101: fc_kernel = 8'h04;
     14'b00100110110110: fc_kernel = 8'h07;
     14'b00100110110111: fc_kernel = 8'h03;
     14'b00100110111000: fc_kernel = 8'h07;
     14'b00100110111001: fc_kernel = 8'h06;
     14'b00100110111010: fc_kernel = 8'h05;
     14'b00100110111011: fc_kernel = 8'h08;
     14'b00100110111100: fc_kernel = 8'h04;
     14'b00100110111101: fc_kernel = 8'h03;
     14'b00100110111110: fc_kernel = 8'h06;
     14'b00100110111111: fc_kernel = 8'h02;
     14'b00100111000000: fc_kernel = 8'h00;
     14'b00100111000001: fc_kernel = 8'h04;
     14'b00100111000010: fc_kernel = 8'h07;
     14'b00100111000011: fc_kernel = 8'h09;
     14'b00100111000100: fc_kernel = 8'h0f;
     14'b00100111000101: fc_kernel = 8'h0c;
     14'b00100111000110: fc_kernel = 8'h0b;
     14'b00100111000111: fc_kernel = 8'h22;
     14'b00100111001000: fc_kernel = 8'h05;
     14'b00100111001001: fc_kernel = 8'h05;
     14'b00100111001010: fc_kernel = 8'h00;
     14'b00100111001011: fc_kernel = 8'h05;
     14'b00100111001100: fc_kernel = 8'h04;
     14'b00100111001101: fc_kernel = 8'h04;
     14'b00100111001110: fc_kernel = 8'h0a;
     14'b00100111001111: fc_kernel = 8'h05;
     14'b00100111010000: fc_kernel = 8'h0a;
     14'b00100111010001: fc_kernel = 8'h0b;
     14'b00100111010010: fc_kernel = 8'h09;
     14'b00100111010011: fc_kernel = 8'h03;
     14'b00100111010100: fc_kernel = 8'hfd;
     14'b00100111010101: fc_kernel = 8'hfe;
     14'b00100111010110: fc_kernel = 8'h03;
     14'b00100111010111: fc_kernel = 8'h04;
     14'b00100111011000: fc_kernel = 8'h09;
     14'b00100111011001: fc_kernel = 8'h09;
     14'b00100111011010: fc_kernel = 8'h05;
     14'b00100111011011: fc_kernel = 8'h03;
     14'b00100111011100: fc_kernel = 8'h07;
     14'b00100111011101: fc_kernel = 8'h04;
     14'b00100111011110: fc_kernel = 8'h0e;
     14'b00100111011111: fc_kernel = 8'h15;
     14'b00100111100000: fc_kernel = 8'h13;
     14'b00100111100001: fc_kernel = 8'h0b;
     14'b00100111100010: fc_kernel = 8'h06;
     14'b00100111100011: fc_kernel = 8'h0c;
     14'b00100111100100: fc_kernel = 8'h08;
     14'b00100111100101: fc_kernel = 8'h07;
     14'b00100111100110: fc_kernel = 8'h09;
     14'b00100111100111: fc_kernel = 8'h07;
     14'b00100111101000: fc_kernel = 8'h07;
     14'b00100111101001: fc_kernel = 8'h09;
     14'b00100111101010: fc_kernel = 8'h02;
     14'b00100111101011: fc_kernel = 8'hfe;
     14'b00100111101100: fc_kernel = 8'hfd;
     14'b00100111101101: fc_kernel = 8'hfd;
     14'b00100111101110: fc_kernel = 8'hff;
     14'b00100111101111: fc_kernel = 8'h06;
     14'b00100111110000: fc_kernel = 8'h05;
     14'b00100111110001: fc_kernel = 8'h0d;
     14'b00100111110010: fc_kernel = 8'h09;
     14'b00100111110011: fc_kernel = 8'h05;
     14'b00100111110100: fc_kernel = 8'h0e;
     14'b00100111110101: fc_kernel = 8'h0b;
     14'b00100111110110: fc_kernel = 8'h0c;
     14'b00100111110111: fc_kernel = 8'h0d;
     14'b00100111111000: fc_kernel = 8'h04;
     14'b00100111111001: fc_kernel = 8'h08;
     14'b00100111111010: fc_kernel = 8'hfe;
     14'b00100111111011: fc_kernel = 8'hff;
     14'b00100111111100: fc_kernel = 8'h03;
     14'b00100111111101: fc_kernel = 8'h08;
     14'b00100111111110: fc_kernel = 8'h0c;
     14'b00100111111111: fc_kernel = 8'h0e;
     14'b00101000000000: fc_kernel = 8'h08;
     14'b00101000000001: fc_kernel = 8'h09;
     14'b00101000000010: fc_kernel = 8'h08;
     14'b00101000000011: fc_kernel = 8'h01;
     14'b00101000000100: fc_kernel = 8'h02;
     14'b00101000000101: fc_kernel = 8'hfc;
     14'b00101000000110: fc_kernel = 8'hfd;
     14'b00101000000111: fc_kernel = 8'h02;
     14'b00101000001000: fc_kernel = 8'h09;
     14'b00101000001001: fc_kernel = 8'h0e;
     14'b00101000001010: fc_kernel = 8'h0c;
     14'b00101000001011: fc_kernel = 8'h14;
     14'b00101000001100: fc_kernel = 8'h0e;
     14'b00101000001101: fc_kernel = 8'h12;
     14'b00101000001110: fc_kernel = 8'h11;
     14'b00101000001111: fc_kernel = 8'h15;
     14'b00101000010000: fc_kernel = 8'h02;
     14'b00101000010001: fc_kernel = 8'hfc;
     14'b00101000010010: fc_kernel = 8'hf6;
     14'b00101000010011: fc_kernel = 8'hfa;
     14'b00101000010100: fc_kernel = 8'hfa;
     14'b00101000010101: fc_kernel = 8'hff;
     14'b00101000010110: fc_kernel = 8'hff;
     14'b00101000010111: fc_kernel = 8'h00;
     14'b00101000011000: fc_kernel = 8'hfa;
     14'b00101000011001: fc_kernel = 8'hfd;
     14'b00101000011010: fc_kernel = 8'h00;
     14'b00101000011011: fc_kernel = 8'h01;
     14'b00101000011100: fc_kernel = 8'h00;
     14'b00101000011101: fc_kernel = 8'h03;
     14'b00101000011110: fc_kernel = 8'h02;
     14'b00101000011111: fc_kernel = 8'h01;
     14'b00101000100000: fc_kernel = 8'h08;
     14'b00101000100001: fc_kernel = 8'h08;
     14'b00101000100010: fc_kernel = 8'h05;
     14'b00101000100011: fc_kernel = 8'h04;
     14'b00101000100100: fc_kernel = 8'h06;
     14'b00101000100101: fc_kernel = 8'h06;
     14'b00101000100110: fc_kernel = 8'h14;
     14'b00101000100111: fc_kernel = 8'h21;
     14'b00101000101000: fc_kernel = 8'hee;
     14'b00101000101001: fc_kernel = 8'hea;
     14'b00101000101010: fc_kernel = 8'he1;
     14'b00101000101011: fc_kernel = 8'hde;
     14'b00101000101100: fc_kernel = 8'he4;
     14'b00101000101101: fc_kernel = 8'he7;
     14'b00101000101110: fc_kernel = 8'he8;
     14'b00101000101111: fc_kernel = 8'he8;
     14'b00101000110000: fc_kernel = 8'hee;
     14'b00101000110001: fc_kernel = 8'heb;
     14'b00101000110010: fc_kernel = 8'hef;
     14'b00101000110011: fc_kernel = 8'hf8;
     14'b00101000110100: fc_kernel = 8'hfb;
     14'b00101000110101: fc_kernel = 8'h00;
     14'b00101000110110: fc_kernel = 8'hfe;
     14'b00101000110111: fc_kernel = 8'h00;
     14'b00101000111000: fc_kernel = 8'hf9;
     14'b00101000111001: fc_kernel = 8'hf3;
     14'b00101000111010: fc_kernel = 8'hf5;
     14'b00101000111011: fc_kernel = 8'hf5;
     14'b00101000111100: fc_kernel = 8'hf3;
     14'b00101000111101: fc_kernel = 8'hf6;
     14'b00101000111110: fc_kernel = 8'h0f;
     14'b00101000111111: fc_kernel = 8'h24;
     14'b00110000000000: fc_kernel = 8'h02;
     14'b00110000000001: fc_kernel = 8'h13;
     14'b00110000000010: fc_kernel = 8'h04;
     14'b00110000000011: fc_kernel = 8'h13;
     14'b00110000000100: fc_kernel = 8'h04;
     14'b00110000000101: fc_kernel = 8'hef;
     14'b00110000000110: fc_kernel = 8'h0f;
     14'b00110000000111: fc_kernel = 8'hff;
     14'b00110000001000: fc_kernel = 8'h09;
     14'b00110000001001: fc_kernel = 8'h10;
     14'b00110000001010: fc_kernel = 8'h13;
     14'b00110000001011: fc_kernel = 8'h0d;
     14'b00110000001100: fc_kernel = 8'h01;
     14'b00110000001101: fc_kernel = 8'hf9;
     14'b00110000001110: fc_kernel = 8'h02;
     14'b00110000001111: fc_kernel = 8'hfc;
     14'b00110000010000: fc_kernel = 8'hf2;
     14'b00110000010001: fc_kernel = 8'hef;
     14'b00110000010010: fc_kernel = 8'hee;
     14'b00110000010011: fc_kernel = 8'hf1;
     14'b00110000010100: fc_kernel = 8'hea;
     14'b00110000010101: fc_kernel = 8'he6;
     14'b00110000010110: fc_kernel = 8'he8;
     14'b00110000010111: fc_kernel = 8'hda;
     14'b00110000011000: fc_kernel = 8'h0c;
     14'b00110000011001: fc_kernel = 8'h03;
     14'b00110000011010: fc_kernel = 8'h11;
     14'b00110000011011: fc_kernel = 8'h11;
     14'b00110000011100: fc_kernel = 8'h08;
     14'b00110000011101: fc_kernel = 8'h17;
     14'b00110000011110: fc_kernel = 8'h13;
     14'b00110000011111: fc_kernel = 8'h0c;
     14'b00110000100000: fc_kernel = 8'h0a;
     14'b00110000100001: fc_kernel = 8'h16;
     14'b00110000100010: fc_kernel = 8'h12;
     14'b00110000100011: fc_kernel = 8'h17;
     14'b00110000100100: fc_kernel = 8'h10;
     14'b00110000100101: fc_kernel = 8'h0b;
     14'b00110000100110: fc_kernel = 8'h08;
     14'b00110000100111: fc_kernel = 8'h0a;
     14'b00110000101000: fc_kernel = 8'h02;
     14'b00110000101001: fc_kernel = 8'h04;
     14'b00110000101010: fc_kernel = 8'h02;
     14'b00110000101011: fc_kernel = 8'hed;
     14'b00110000101100: fc_kernel = 8'hd7;
     14'b00110000101101: fc_kernel = 8'hcf;
     14'b00110000101110: fc_kernel = 8'hdf;
     14'b00110000101111: fc_kernel = 8'he2;
     14'b00110000110000: fc_kernel = 8'hff;
     14'b00110000110001: fc_kernel = 8'h11;
     14'b00110000110010: fc_kernel = 8'h18;
     14'b00110000110011: fc_kernel = 8'h17;
     14'b00110000110100: fc_kernel = 8'h14;
     14'b00110000110101: fc_kernel = 8'h0f;
     14'b00110000110110: fc_kernel = 8'h08;
     14'b00110000110111: fc_kernel = 8'h0a;
     14'b00110000111000: fc_kernel = 8'h09;
     14'b00110000111001: fc_kernel = 8'h11;
     14'b00110000111010: fc_kernel = 8'h0c;
     14'b00110000111011: fc_kernel = 8'h0e;
     14'b00110000111100: fc_kernel = 8'h09;
     14'b00110000111101: fc_kernel = 8'h09;
     14'b00110000111110: fc_kernel = 8'h0a;
     14'b00110000111111: fc_kernel = 8'h00;
     14'b00110001000000: fc_kernel = 8'h03;
     14'b00110001000001: fc_kernel = 8'h06;
     14'b00110001000010: fc_kernel = 8'h00;
     14'b00110001000011: fc_kernel = 8'hfc;
     14'b00110001000100: fc_kernel = 8'hee;
     14'b00110001000101: fc_kernel = 8'hd8;
     14'b00110001000110: fc_kernel = 8'hc3;
     14'b00110001000111: fc_kernel = 8'hda;
     14'b00110001001000: fc_kernel = 8'h1a;
     14'b00110001001001: fc_kernel = 8'h12;
     14'b00110001001010: fc_kernel = 8'h11;
     14'b00110001001011: fc_kernel = 8'h11;
     14'b00110001001100: fc_kernel = 8'h0e;
     14'b00110001001101: fc_kernel = 8'h09;
     14'b00110001001110: fc_kernel = 8'h07;
     14'b00110001001111: fc_kernel = 8'h0b;
     14'b00110001010000: fc_kernel = 8'h0e;
     14'b00110001010001: fc_kernel = 8'h07;
     14'b00110001010010: fc_kernel = 8'h07;
     14'b00110001010011: fc_kernel = 8'h06;
     14'b00110001010100: fc_kernel = 8'h00;
     14'b00110001010101: fc_kernel = 8'h04;
     14'b00110001010110: fc_kernel = 8'h03;
     14'b00110001010111: fc_kernel = 8'hff;
     14'b00110001011000: fc_kernel = 8'h01;
     14'b00110001011001: fc_kernel = 8'h01;
     14'b00110001011010: fc_kernel = 8'hfc;
     14'b00110001011011: fc_kernel = 8'hf9;
     14'b00110001011100: fc_kernel = 8'hf2;
     14'b00110001011101: fc_kernel = 8'hf3;
     14'b00110001011110: fc_kernel = 8'hdc;
     14'b00110001011111: fc_kernel = 8'hcc;
     14'b00110001100000: fc_kernel = 8'h11;
     14'b00110001100001: fc_kernel = 8'h06;
     14'b00110001100010: fc_kernel = 8'h12;
     14'b00110001100011: fc_kernel = 8'h11;
     14'b00110001100100: fc_kernel = 8'h08;
     14'b00110001100101: fc_kernel = 8'h09;
     14'b00110001100110: fc_kernel = 8'h05;
     14'b00110001100111: fc_kernel = 8'h07;
     14'b00110001101000: fc_kernel = 8'h09;
     14'b00110001101001: fc_kernel = 8'h02;
     14'b00110001101010: fc_kernel = 8'h03;
     14'b00110001101011: fc_kernel = 8'h03;
     14'b00110001101100: fc_kernel = 8'h07;
     14'b00110001101101: fc_kernel = 8'h08;
     14'b00110001101110: fc_kernel = 8'h07;
     14'b00110001101111: fc_kernel = 8'h06;
     14'b00110001110000: fc_kernel = 8'h00;
     14'b00110001110001: fc_kernel = 8'hfd;
     14'b00110001110010: fc_kernel = 8'hfa;
     14'b00110001110011: fc_kernel = 8'hf7;
     14'b00110001110100: fc_kernel = 8'hf8;
     14'b00110001110101: fc_kernel = 8'hf2;
     14'b00110001110110: fc_kernel = 8'hee;
     14'b00110001110111: fc_kernel = 8'he9;
     14'b00110001111000: fc_kernel = 8'h0f;
     14'b00110001111001: fc_kernel = 8'h04;
     14'b00110001111010: fc_kernel = 8'h10;
     14'b00110001111011: fc_kernel = 8'h0a;
     14'b00110001111100: fc_kernel = 8'h08;
     14'b00110001111101: fc_kernel = 8'h05;
     14'b00110001111110: fc_kernel = 8'h00;
     14'b00110001111111: fc_kernel = 8'h03;
     14'b00110010000000: fc_kernel = 8'h06;
     14'b00110010000001: fc_kernel = 8'h02;
     14'b00110010000010: fc_kernel = 8'h04;
     14'b00110010000011: fc_kernel = 8'h08;
     14'b00110010000100: fc_kernel = 8'h07;
     14'b00110010000101: fc_kernel = 8'h05;
     14'b00110010000110: fc_kernel = 8'h02;
     14'b00110010000111: fc_kernel = 8'h00;
     14'b00110010001000: fc_kernel = 8'h03;
     14'b00110010001001: fc_kernel = 8'hff;
     14'b00110010001010: fc_kernel = 8'hff;
     14'b00110010001011: fc_kernel = 8'hf9;
     14'b00110010001100: fc_kernel = 8'hf2;
     14'b00110010001101: fc_kernel = 8'hf3;
     14'b00110010001110: fc_kernel = 8'hea;
     14'b00110010001111: fc_kernel = 8'he7;
     14'b00110010010000: fc_kernel = 8'h01;
     14'b00110010010001: fc_kernel = 8'h09;
     14'b00110010010010: fc_kernel = 8'h0f;
     14'b00110010010011: fc_kernel = 8'h0c;
     14'b00110010010100: fc_kernel = 8'h04;
     14'b00110010010101: fc_kernel = 8'h00;
     14'b00110010010110: fc_kernel = 8'h01;
     14'b00110010010111: fc_kernel = 8'h00;
     14'b00110010011000: fc_kernel = 8'h04;
     14'b00110010011001: fc_kernel = 8'h07;
     14'b00110010011010: fc_kernel = 8'h06;
     14'b00110010011011: fc_kernel = 8'h09;
     14'b00110010011100: fc_kernel = 8'h07;
     14'b00110010011101: fc_kernel = 8'h0b;
     14'b00110010011110: fc_kernel = 8'h01;
     14'b00110010011111: fc_kernel = 8'h07;
     14'b00110010100000: fc_kernel = 8'h00;
     14'b00110010100001: fc_kernel = 8'h07;
     14'b00110010100010: fc_kernel = 8'h00;
     14'b00110010100011: fc_kernel = 8'h03;
     14'b00110010100100: fc_kernel = 8'hfb;
     14'b00110010100101: fc_kernel = 8'hed;
     14'b00110010100110: fc_kernel = 8'hd6;
     14'b00110010100111: fc_kernel = 8'hc6;
     14'b00110010101000: fc_kernel = 8'h0c;
     14'b00110010101001: fc_kernel = 8'h0e;
     14'b00110010101010: fc_kernel = 8'h0e;
     14'b00110010101011: fc_kernel = 8'h02;
     14'b00110010101100: fc_kernel = 8'h04;
     14'b00110010101101: fc_kernel = 8'h08;
     14'b00110010101110: fc_kernel = 8'h05;
     14'b00110010101111: fc_kernel = 8'h00;
     14'b00110010110000: fc_kernel = 8'h00;
     14'b00110010110001: fc_kernel = 8'hfd;
     14'b00110010110010: fc_kernel = 8'hfa;
     14'b00110010110011: fc_kernel = 8'h01;
     14'b00110010110100: fc_kernel = 8'h07;
     14'b00110010110101: fc_kernel = 8'h0b;
     14'b00110010110110: fc_kernel = 8'h05;
     14'b00110010110111: fc_kernel = 8'h05;
     14'b00110010111000: fc_kernel = 8'h05;
     14'b00110010111001: fc_kernel = 8'h04;
     14'b00110010111010: fc_kernel = 8'h04;
     14'b00110010111011: fc_kernel = 8'h04;
     14'b00110010111100: fc_kernel = 8'h05;
     14'b00110010111101: fc_kernel = 8'hfa;
     14'b00110010111110: fc_kernel = 8'hcd;
     14'b00110010111111: fc_kernel = 8'ha9;
     14'b00110011000000: fc_kernel = 8'h14;
     14'b00110011000001: fc_kernel = 8'h16;
     14'b00110011000010: fc_kernel = 8'h0c;
     14'b00110011000011: fc_kernel = 8'h01;
     14'b00110011000100: fc_kernel = 8'h02;
     14'b00110011000101: fc_kernel = 8'h00;
     14'b00110011000110: fc_kernel = 8'hfc;
     14'b00110011000111: fc_kernel = 8'hf9;
     14'b00110011001000: fc_kernel = 8'hf1;
     14'b00110011001001: fc_kernel = 8'hf1;
     14'b00110011001010: fc_kernel = 8'hf2;
     14'b00110011001011: fc_kernel = 8'hf8;
     14'b00110011001100: fc_kernel = 8'h05;
     14'b00110011001101: fc_kernel = 8'h0a;
     14'b00110011001110: fc_kernel = 8'h05;
     14'b00110011001111: fc_kernel = 8'h07;
     14'b00110011010000: fc_kernel = 8'h05;
     14'b00110011010001: fc_kernel = 8'h08;
     14'b00110011010010: fc_kernel = 8'h08;
     14'b00110011010011: fc_kernel = 8'h08;
     14'b00110011010100: fc_kernel = 8'h08;
     14'b00110011010101: fc_kernel = 8'h03;
     14'b00110011010110: fc_kernel = 8'he0;
     14'b00110011010111: fc_kernel = 8'hb3;
     14'b00110011011000: fc_kernel = 8'h1a;
     14'b00110011011001: fc_kernel = 8'h21;
     14'b00110011011010: fc_kernel = 8'h0b;
     14'b00110011011011: fc_kernel = 8'h02;
     14'b00110011011100: fc_kernel = 8'hfb;
     14'b00110011011101: fc_kernel = 8'hf4;
     14'b00110011011110: fc_kernel = 8'hed;
     14'b00110011011111: fc_kernel = 8'heb;
     14'b00110011100000: fc_kernel = 8'hee;
     14'b00110011100001: fc_kernel = 8'hf0;
     14'b00110011100010: fc_kernel = 8'hf5;
     14'b00110011100011: fc_kernel = 8'h01;
     14'b00110011100100: fc_kernel = 8'h0f;
     14'b00110011100101: fc_kernel = 8'h05;
     14'b00110011100110: fc_kernel = 8'h08;
     14'b00110011100111: fc_kernel = 8'h05;
     14'b00110011101000: fc_kernel = 8'h06;
     14'b00110011101001: fc_kernel = 8'h06;
     14'b00110011101010: fc_kernel = 8'h05;
     14'b00110011101011: fc_kernel = 8'h04;
     14'b00110011101100: fc_kernel = 8'h07;
     14'b00110011101101: fc_kernel = 8'h01;
     14'b00110011101110: fc_kernel = 8'he8;
     14'b00110011101111: fc_kernel = 8'hce;
     14'b00110011110000: fc_kernel = 8'h10;
     14'b00110011110001: fc_kernel = 8'h0f;
     14'b00110011110010: fc_kernel = 8'h00;
     14'b00110011110011: fc_kernel = 8'hfe;
     14'b00110011110100: fc_kernel = 8'hf6;
     14'b00110011110101: fc_kernel = 8'hf0;
     14'b00110011110110: fc_kernel = 8'hf0;
     14'b00110011110111: fc_kernel = 8'hf3;
     14'b00110011111000: fc_kernel = 8'hfa;
     14'b00110011111001: fc_kernel = 8'hfd;
     14'b00110011111010: fc_kernel = 8'hff;
     14'b00110011111011: fc_kernel = 8'h09;
     14'b00110011111100: fc_kernel = 8'h0c;
     14'b00110011111101: fc_kernel = 8'h02;
     14'b00110011111110: fc_kernel = 8'h07;
     14'b00110011111111: fc_kernel = 8'h02;
     14'b00110100000000: fc_kernel = 8'h03;
     14'b00110100000001: fc_kernel = 8'h04;
     14'b00110100000010: fc_kernel = 8'hfc;
     14'b00110100000011: fc_kernel = 8'hf6;
     14'b00110100000100: fc_kernel = 8'hee;
     14'b00110100000101: fc_kernel = 8'hf0;
     14'b00110100000110: fc_kernel = 8'he9;
     14'b00110100000111: fc_kernel = 8'he5;
     14'b00110100001000: fc_kernel = 8'h0d;
     14'b00110100001001: fc_kernel = 8'h05;
     14'b00110100001010: fc_kernel = 8'hf7;
     14'b00110100001011: fc_kernel = 8'hf4;
     14'b00110100001100: fc_kernel = 8'heb;
     14'b00110100001101: fc_kernel = 8'hf2;
     14'b00110100001110: fc_kernel = 8'hf7;
     14'b00110100001111: fc_kernel = 8'hfa;
     14'b00110100010000: fc_kernel = 8'hfa;
     14'b00110100010001: fc_kernel = 8'hfa;
     14'b00110100010010: fc_kernel = 8'h01;
     14'b00110100010011: fc_kernel = 8'h09;
     14'b00110100010100: fc_kernel = 8'h08;
     14'b00110100010101: fc_kernel = 8'hfe;
     14'b00110100010110: fc_kernel = 8'h00;
     14'b00110100010111: fc_kernel = 8'h07;
     14'b00110100011000: fc_kernel = 8'h03;
     14'b00110100011001: fc_kernel = 8'h01;
     14'b00110100011010: fc_kernel = 8'hf6;
     14'b00110100011011: fc_kernel = 8'he6;
     14'b00110100011100: fc_kernel = 8'hdb;
     14'b00110100011101: fc_kernel = 8'hdd;
     14'b00110100011110: fc_kernel = 8'he7;
     14'b00110100011111: fc_kernel = 8'heb;
     14'b00110100100000: fc_kernel = 8'h11;
     14'b00110100100001: fc_kernel = 8'hfc;
     14'b00110100100010: fc_kernel = 8'hf9;
     14'b00110100100011: fc_kernel = 8'hf3;
     14'b00110100100100: fc_kernel = 8'hf1;
     14'b00110100100101: fc_kernel = 8'hf1;
     14'b00110100100110: fc_kernel = 8'hf9;
     14'b00110100100111: fc_kernel = 8'hf9;
     14'b00110100101000: fc_kernel = 8'hf8;
     14'b00110100101001: fc_kernel = 8'hf4;
     14'b00110100101010: fc_kernel = 8'hfc;
     14'b00110100101011: fc_kernel = 8'h05;
     14'b00110100101100: fc_kernel = 8'h04;
     14'b00110100101101: fc_kernel = 8'h03;
     14'b00110100101110: fc_kernel = 8'h03;
     14'b00110100101111: fc_kernel = 8'h01;
     14'b00110100110000: fc_kernel = 8'h04;
     14'b00110100110001: fc_kernel = 8'hfb;
     14'b00110100110010: fc_kernel = 8'hf4;
     14'b00110100110011: fc_kernel = 8'hf3;
     14'b00110100110100: fc_kernel = 8'hed;
     14'b00110100110101: fc_kernel = 8'he7;
     14'b00110100110110: fc_kernel = 8'hf0;
     14'b00110100110111: fc_kernel = 8'hef;
     14'b00110100111000: fc_kernel = 8'h10;
     14'b00110100111001: fc_kernel = 8'h00;
     14'b00110100111010: fc_kernel = 8'hfc;
     14'b00110100111011: fc_kernel = 8'hf0;
     14'b00110100111100: fc_kernel = 8'hed;
     14'b00110100111101: fc_kernel = 8'hee;
     14'b00110100111110: fc_kernel = 8'hf3;
     14'b00110100111111: fc_kernel = 8'hf8;
     14'b00110101000000: fc_kernel = 8'hfb;
     14'b00110101000001: fc_kernel = 8'hfc;
     14'b00110101000010: fc_kernel = 8'h02;
     14'b00110101000011: fc_kernel = 8'h0a;
     14'b00110101000100: fc_kernel = 8'h01;
     14'b00110101000101: fc_kernel = 8'h01;
     14'b00110101000110: fc_kernel = 8'hfd;
     14'b00110101000111: fc_kernel = 8'h01;
     14'b00110101001000: fc_kernel = 8'hfe;
     14'b00110101001001: fc_kernel = 8'hfe;
     14'b00110101001010: fc_kernel = 8'h01;
     14'b00110101001011: fc_kernel = 8'hff;
     14'b00110101001100: fc_kernel = 8'hfa;
     14'b00110101001101: fc_kernel = 8'h01;
     14'b00110101001110: fc_kernel = 8'h03;
     14'b00110101001111: fc_kernel = 8'hf3;
     14'b00110101010000: fc_kernel = 8'h0c;
     14'b00110101010001: fc_kernel = 8'h0f;
     14'b00110101010010: fc_kernel = 8'h03;
     14'b00110101010011: fc_kernel = 8'h00;
     14'b00110101010100: fc_kernel = 8'hf7;
     14'b00110101010101: fc_kernel = 8'hf0;
     14'b00110101010110: fc_kernel = 8'hef;
     14'b00110101010111: fc_kernel = 8'hf6;
     14'b00110101011000: fc_kernel = 8'hf6;
     14'b00110101011001: fc_kernel = 8'h00;
     14'b00110101011010: fc_kernel = 8'h03;
     14'b00110101011011: fc_kernel = 8'h03;
     14'b00110101011100: fc_kernel = 8'h00;
     14'b00110101011101: fc_kernel = 8'hfc;
     14'b00110101011110: fc_kernel = 8'hf6;
     14'b00110101011111: fc_kernel = 8'hfe;
     14'b00110101100000: fc_kernel = 8'hfd;
     14'b00110101100001: fc_kernel = 8'h00;
     14'b00110101100010: fc_kernel = 8'h01;
     14'b00110101100011: fc_kernel = 8'hfc;
     14'b00110101100100: fc_kernel = 8'hfc;
     14'b00110101100101: fc_kernel = 8'h0a;
     14'b00110101100110: fc_kernel = 8'h15;
     14'b00110101100111: fc_kernel = 8'hf8;
     14'b00110101101000: fc_kernel = 8'h11;
     14'b00110101101001: fc_kernel = 8'h18;
     14'b00110101101010: fc_kernel = 8'h0e;
     14'b00110101101011: fc_kernel = 8'h03;
     14'b00110101101100: fc_kernel = 8'hfb;
     14'b00110101101101: fc_kernel = 8'hf5;
     14'b00110101101110: fc_kernel = 8'hf1;
     14'b00110101101111: fc_kernel = 8'he7;
     14'b00110101110000: fc_kernel = 8'hed;
     14'b00110101110001: fc_kernel = 8'hf3;
     14'b00110101110010: fc_kernel = 8'hfc;
     14'b00110101110011: fc_kernel = 8'hfd;
     14'b00110101110100: fc_kernel = 8'hf9;
     14'b00110101110101: fc_kernel = 8'hf2;
     14'b00110101110110: fc_kernel = 8'hfb;
     14'b00110101110111: fc_kernel = 8'hfb;
     14'b00110101111000: fc_kernel = 8'h02;
     14'b00110101111001: fc_kernel = 8'h04;
     14'b00110101111010: fc_kernel = 8'h00;
     14'b00110101111011: fc_kernel = 8'hfc;
     14'b00110101111100: fc_kernel = 8'h06;
     14'b00110101111101: fc_kernel = 8'h09;
     14'b00110101111110: fc_kernel = 8'hfd;
     14'b00110101111111: fc_kernel = 8'he3;
     14'b00110110000000: fc_kernel = 8'h1f;
     14'b00110110000001: fc_kernel = 8'h19;
     14'b00110110000010: fc_kernel = 8'h11;
     14'b00110110000011: fc_kernel = 8'h08;
     14'b00110110000100: fc_kernel = 8'hfd;
     14'b00110110000101: fc_kernel = 8'hfb;
     14'b00110110000110: fc_kernel = 8'hf2;
     14'b00110110000111: fc_kernel = 8'hec;
     14'b00110110001000: fc_kernel = 8'he7;
     14'b00110110001001: fc_kernel = 8'hed;
     14'b00110110001010: fc_kernel = 8'hee;
     14'b00110110001011: fc_kernel = 8'hf3;
     14'b00110110001100: fc_kernel = 8'hf0;
     14'b00110110001101: fc_kernel = 8'hfa;
     14'b00110110001110: fc_kernel = 8'h04;
     14'b00110110001111: fc_kernel = 8'h04;
     14'b00110110010000: fc_kernel = 8'h05;
     14'b00110110010001: fc_kernel = 8'hfd;
     14'b00110110010010: fc_kernel = 8'hff;
     14'b00110110010011: fc_kernel = 8'hff;
     14'b00110110010100: fc_kernel = 8'h06;
     14'b00110110010101: fc_kernel = 8'h06;
     14'b00110110010110: fc_kernel = 8'hf6;
     14'b00110110010111: fc_kernel = 8'hd2;
     14'b00110110011000: fc_kernel = 8'h16;
     14'b00110110011001: fc_kernel = 8'h12;
     14'b00110110011010: fc_kernel = 8'h12;
     14'b00110110011011: fc_kernel = 8'h0b;
     14'b00110110011100: fc_kernel = 8'h02;
     14'b00110110011101: fc_kernel = 8'h00;
     14'b00110110011110: fc_kernel = 8'hfc;
     14'b00110110011111: fc_kernel = 8'hf5;
     14'b00110110100000: fc_kernel = 8'hef;
     14'b00110110100001: fc_kernel = 8'hf0;
     14'b00110110100010: fc_kernel = 8'he9;
     14'b00110110100011: fc_kernel = 8'hf2;
     14'b00110110100100: fc_kernel = 8'hf9;
     14'b00110110100101: fc_kernel = 8'h00;
     14'b00110110100110: fc_kernel = 8'h08;
     14'b00110110100111: fc_kernel = 8'h09;
     14'b00110110101000: fc_kernel = 8'h05;
     14'b00110110101001: fc_kernel = 8'h01;
     14'b00110110101010: fc_kernel = 8'h00;
     14'b00110110101011: fc_kernel = 8'h05;
     14'b00110110101100: fc_kernel = 8'h04;
     14'b00110110101101: fc_kernel = 8'h00;
     14'b00110110101110: fc_kernel = 8'hf9;
     14'b00110110101111: fc_kernel = 8'he3;
     14'b00110110110000: fc_kernel = 8'h0a;
     14'b00110110110001: fc_kernel = 8'h0d;
     14'b00110110110010: fc_kernel = 8'h0b;
     14'b00110110110011: fc_kernel = 8'h07;
     14'b00110110110100: fc_kernel = 8'h0e;
     14'b00110110110101: fc_kernel = 8'h01;
     14'b00110110110110: fc_kernel = 8'h03;
     14'b00110110110111: fc_kernel = 8'h05;
     14'b00110110111000: fc_kernel = 8'hfd;
     14'b00110110111001: fc_kernel = 8'hf3;
     14'b00110110111010: fc_kernel = 8'hf3;
     14'b00110110111011: fc_kernel = 8'hf9;
     14'b00110110111100: fc_kernel = 8'h00;
     14'b00110110111101: fc_kernel = 8'hfe;
     14'b00110110111110: fc_kernel = 8'h04;
     14'b00110110111111: fc_kernel = 8'h03;
     14'b00110111000000: fc_kernel = 8'h07;
     14'b00110111000001: fc_kernel = 8'h05;
     14'b00110111000010: fc_kernel = 8'h01;
     14'b00110111000011: fc_kernel = 8'h00;
     14'b00110111000100: fc_kernel = 8'hfa;
     14'b00110111000101: fc_kernel = 8'hfe;
     14'b00110111000110: fc_kernel = 8'hf6;
     14'b00110111000111: fc_kernel = 8'he3;
     14'b00110111001000: fc_kernel = 8'h0c;
     14'b00110111001001: fc_kernel = 8'h09;
     14'b00110111001010: fc_kernel = 8'h0e;
     14'b00110111001011: fc_kernel = 8'h03;
     14'b00110111001100: fc_kernel = 8'h04;
     14'b00110111001101: fc_kernel = 8'h08;
     14'b00110111001110: fc_kernel = 8'hfe;
     14'b00110111001111: fc_kernel = 8'h00;
     14'b00110111010000: fc_kernel = 8'hf8;
     14'b00110111010001: fc_kernel = 8'hfa;
     14'b00110111010010: fc_kernel = 8'hf6;
     14'b00110111010011: fc_kernel = 8'hf6;
     14'b00110111010100: fc_kernel = 8'hff;
     14'b00110111010101: fc_kernel = 8'h00;
     14'b00110111010110: fc_kernel = 8'h06;
     14'b00110111010111: fc_kernel = 8'h05;
     14'b00110111011000: fc_kernel = 8'h08;
     14'b00110111011001: fc_kernel = 8'h02;
     14'b00110111011010: fc_kernel = 8'h03;
     14'b00110111011011: fc_kernel = 8'hff;
     14'b00110111011100: fc_kernel = 8'hf8;
     14'b00110111011101: fc_kernel = 8'hfb;
     14'b00110111011110: fc_kernel = 8'hee;
     14'b00110111011111: fc_kernel = 8'he2;
     14'b00110111100000: fc_kernel = 8'h12;
     14'b00110111100001: fc_kernel = 8'h0f;
     14'b00110111100010: fc_kernel = 8'h08;
     14'b00110111100011: fc_kernel = 8'h04;
     14'b00110111100100: fc_kernel = 8'h06;
     14'b00110111100101: fc_kernel = 8'h06;
     14'b00110111100110: fc_kernel = 8'h04;
     14'b00110111100111: fc_kernel = 8'h02;
     14'b00110111101000: fc_kernel = 8'hfe;
     14'b00110111101001: fc_kernel = 8'hff;
     14'b00110111101010: fc_kernel = 8'hfe;
     14'b00110111101011: fc_kernel = 8'hf9;
     14'b00110111101100: fc_kernel = 8'hfa;
     14'b00110111101101: fc_kernel = 8'h03;
     14'b00110111101110: fc_kernel = 8'h00;
     14'b00110111101111: fc_kernel = 8'h04;
     14'b00110111110000: fc_kernel = 8'h07;
     14'b00110111110001: fc_kernel = 8'h05;
     14'b00110111110010: fc_kernel = 8'h03;
     14'b00110111110011: fc_kernel = 8'hfc;
     14'b00110111110100: fc_kernel = 8'hfc;
     14'b00110111110101: fc_kernel = 8'hf4;
     14'b00110111110110: fc_kernel = 8'he3;
     14'b00110111110111: fc_kernel = 8'hd8;
     14'b00110111111000: fc_kernel = 8'h23;
     14'b00110111111001: fc_kernel = 8'h1f;
     14'b00110111111010: fc_kernel = 8'h11;
     14'b00110111111011: fc_kernel = 8'h08;
     14'b00110111111100: fc_kernel = 8'h09;
     14'b00110111111101: fc_kernel = 8'h05;
     14'b00110111111110: fc_kernel = 8'hfa;
     14'b00110111111111: fc_kernel = 8'hff;
     14'b00111000000000: fc_kernel = 8'hff;
     14'b00111000000001: fc_kernel = 8'h00;
     14'b00111000000010: fc_kernel = 8'hf8;
     14'b00111000000011: fc_kernel = 8'hfd;
     14'b00111000000100: fc_kernel = 8'h02;
     14'b00111000000101: fc_kernel = 8'h00;
     14'b00111000000110: fc_kernel = 8'h02;
     14'b00111000000111: fc_kernel = 8'h02;
     14'b00111000001000: fc_kernel = 8'h05;
     14'b00111000001001: fc_kernel = 8'h02;
     14'b00111000001010: fc_kernel = 8'hfd;
     14'b00111000001011: fc_kernel = 8'hfa;
     14'b00111000001100: fc_kernel = 8'hf5;
     14'b00111000001101: fc_kernel = 8'hf6;
     14'b00111000001110: fc_kernel = 8'he5;
     14'b00111000001111: fc_kernel = 8'hde;
     14'b00111000010000: fc_kernel = 8'h16;
     14'b00111000010001: fc_kernel = 8'h17;
     14'b00111000010010: fc_kernel = 8'h0f;
     14'b00111000010011: fc_kernel = 8'h0b;
     14'b00111000010100: fc_kernel = 8'h0f;
     14'b00111000010101: fc_kernel = 8'h0e;
     14'b00111000010110: fc_kernel = 8'h0b;
     14'b00111000010111: fc_kernel = 8'h06;
     14'b00111000011000: fc_kernel = 8'h07;
     14'b00111000011001: fc_kernel = 8'h0a;
     14'b00111000011010: fc_kernel = 8'h07;
     14'b00111000011011: fc_kernel = 8'h03;
     14'b00111000011100: fc_kernel = 8'h05;
     14'b00111000011101: fc_kernel = 8'h01;
     14'b00111000011110: fc_kernel = 8'h00;
     14'b00111000011111: fc_kernel = 8'h06;
     14'b00111000100000: fc_kernel = 8'h03;
     14'b00111000100001: fc_kernel = 8'h00;
     14'b00111000100010: fc_kernel = 8'hfd;
     14'b00111000100011: fc_kernel = 8'hf7;
     14'b00111000100100: fc_kernel = 8'hf4;
     14'b00111000100101: fc_kernel = 8'hee;
     14'b00111000100110: fc_kernel = 8'he8;
     14'b00111000100111: fc_kernel = 8'he9;
     14'b00111000101000: fc_kernel = 8'h11;
     14'b00111000101001: fc_kernel = 8'h15;
     14'b00111000101010: fc_kernel = 8'h11;
     14'b00111000101011: fc_kernel = 8'h10;
     14'b00111000101100: fc_kernel = 8'h1d;
     14'b00111000101101: fc_kernel = 8'h20;
     14'b00111000101110: fc_kernel = 8'h1c;
     14'b00111000101111: fc_kernel = 8'h19;
     14'b00111000110000: fc_kernel = 8'h1a;
     14'b00111000110001: fc_kernel = 8'h16;
     14'b00111000110010: fc_kernel = 8'h13;
     14'b00111000110011: fc_kernel = 8'h15;
     14'b00111000110100: fc_kernel = 8'h0e;
     14'b00111000110101: fc_kernel = 8'h09;
     14'b00111000110110: fc_kernel = 8'h08;
     14'b00111000110111: fc_kernel = 8'h0a;
     14'b00111000111000: fc_kernel = 8'hfd;
     14'b00111000111001: fc_kernel = 8'hfa;
     14'b00111000111010: fc_kernel = 8'h00;
     14'b00111000111011: fc_kernel = 8'hf9;
     14'b00111000111100: fc_kernel = 8'hf5;
     14'b00111000111101: fc_kernel = 8'hf8;
     14'b00111000111110: fc_kernel = 8'hee;
     14'b00111000111111: fc_kernel = 8'hf1;
     14'b01000000000000: fc_kernel = 8'hff;
     14'b01000000000001: fc_kernel = 8'he4;
     14'b01000000000010: fc_kernel = 8'he6;
     14'b01000000000011: fc_kernel = 8'hf4;
     14'b01000000000100: fc_kernel = 8'hd1;
     14'b01000000000101: fc_kernel = 8'hd7;
     14'b01000000000110: fc_kernel = 8'hc5;
     14'b01000000000111: fc_kernel = 8'hc8;
     14'b01000000001000: fc_kernel = 8'hc6;
     14'b01000000001001: fc_kernel = 8'hbc;
     14'b01000000001010: fc_kernel = 8'hb0;
     14'b01000000001011: fc_kernel = 8'hd7;
     14'b01000000001100: fc_kernel = 8'he3;
     14'b01000000001101: fc_kernel = 8'hd7;
     14'b01000000001110: fc_kernel = 8'hd6;
     14'b01000000001111: fc_kernel = 8'hd8;
     14'b01000000010000: fc_kernel = 8'hd1;
     14'b01000000010001: fc_kernel = 8'hc5;
     14'b01000000010010: fc_kernel = 8'hd3;
     14'b01000000010011: fc_kernel = 8'he6;
     14'b01000000010100: fc_kernel = 8'he2;
     14'b01000000010101: fc_kernel = 8'he0;
     14'b01000000010110: fc_kernel = 8'he0;
     14'b01000000010111: fc_kernel = 8'hfa;
     14'b01000000011000: fc_kernel = 8'hf8;
     14'b01000000011001: fc_kernel = 8'hf3;
     14'b01000000011010: fc_kernel = 8'hef;
     14'b01000000011011: fc_kernel = 8'hf2;
     14'b01000000011100: fc_kernel = 8'hed;
     14'b01000000011101: fc_kernel = 8'he3;
     14'b01000000011110: fc_kernel = 8'hdd;
     14'b01000000011111: fc_kernel = 8'hd7;
     14'b01000000100000: fc_kernel = 8'hd3;
     14'b01000000100001: fc_kernel = 8'hcd;
     14'b01000000100010: fc_kernel = 8'hcb;
     14'b01000000100011: fc_kernel = 8'hcf;
     14'b01000000100100: fc_kernel = 8'hd7;
     14'b01000000100101: fc_kernel = 8'hdb;
     14'b01000000100110: fc_kernel = 8'he0;
     14'b01000000100111: fc_kernel = 8'he6;
     14'b01000000101000: fc_kernel = 8'hed;
     14'b01000000101001: fc_kernel = 8'hf2;
     14'b01000000101010: fc_kernel = 8'hfa;
     14'b01000000101011: fc_kernel = 8'hfc;
     14'b01000000101100: fc_kernel = 8'hf3;
     14'b01000000101101: fc_kernel = 8'heb;
     14'b01000000101110: fc_kernel = 8'hfe;
     14'b01000000101111: fc_kernel = 8'hff;
     14'b01000000110000: fc_kernel = 8'h01;
     14'b01000000110001: fc_kernel = 8'h00;
     14'b01000000110010: fc_kernel = 8'h03;
     14'b01000000110011: fc_kernel = 8'hf2;
     14'b01000000110100: fc_kernel = 8'hf5;
     14'b01000000110101: fc_kernel = 8'hf8;
     14'b01000000110110: fc_kernel = 8'hf3;
     14'b01000000110111: fc_kernel = 8'he3;
     14'b01000000111000: fc_kernel = 8'he1;
     14'b01000000111001: fc_kernel = 8'hea;
     14'b01000000111010: fc_kernel = 8'hed;
     14'b01000000111011: fc_kernel = 8'heb;
     14'b01000000111100: fc_kernel = 8'hee;
     14'b01000000111101: fc_kernel = 8'hf0;
     14'b01000000111110: fc_kernel = 8'hf0;
     14'b01000000111111: fc_kernel = 8'hf5;
     14'b01000001000000: fc_kernel = 8'hf2;
     14'b01000001000001: fc_kernel = 8'h00;
     14'b01000001000010: fc_kernel = 8'h0f;
     14'b01000001000011: fc_kernel = 8'h15;
     14'b01000001000100: fc_kernel = 8'h16;
     14'b01000001000101: fc_kernel = 8'h1a;
     14'b01000001000110: fc_kernel = 8'h13;
     14'b01000001000111: fc_kernel = 8'h0c;
     14'b01000001001000: fc_kernel = 8'hf1;
     14'b01000001001001: fc_kernel = 8'h0f;
     14'b01000001001010: fc_kernel = 8'h08;
     14'b01000001001011: fc_kernel = 8'hfd;
     14'b01000001001100: fc_kernel = 8'hf1;
     14'b01000001001101: fc_kernel = 8'hf3;
     14'b01000001001110: fc_kernel = 8'hf5;
     14'b01000001001111: fc_kernel = 8'hfa;
     14'b01000001010000: fc_kernel = 8'hf4;
     14'b01000001010001: fc_kernel = 8'hf4;
     14'b01000001010010: fc_kernel = 8'hf1;
     14'b01000001010011: fc_kernel = 8'hf3;
     14'b01000001010100: fc_kernel = 8'hf1;
     14'b01000001010101: fc_kernel = 8'hf4;
     14'b01000001010110: fc_kernel = 8'hf8;
     14'b01000001010111: fc_kernel = 8'hf7;
     14'b01000001011000: fc_kernel = 8'hf8;
     14'b01000001011001: fc_kernel = 8'h00;
     14'b01000001011010: fc_kernel = 8'hfe;
     14'b01000001011011: fc_kernel = 8'hfb;
     14'b01000001011100: fc_kernel = 8'h01;
     14'b01000001011101: fc_kernel = 8'h13;
     14'b01000001011110: fc_kernel = 8'h09;
     14'b01000001011111: fc_kernel = 8'h00;
     14'b01000001100000: fc_kernel = 8'hf2;
     14'b01000001100001: fc_kernel = 8'hf9;
     14'b01000001100010: fc_kernel = 8'h06;
     14'b01000001100011: fc_kernel = 8'h05;
     14'b01000001100100: fc_kernel = 8'hf7;
     14'b01000001100101: fc_kernel = 8'hf6;
     14'b01000001100110: fc_kernel = 8'hfc;
     14'b01000001100111: fc_kernel = 8'hfc;
     14'b01000001101000: fc_kernel = 8'hf4;
     14'b01000001101001: fc_kernel = 8'hf1;
     14'b01000001101010: fc_kernel = 8'heb;
     14'b01000001101011: fc_kernel = 8'hef;
     14'b01000001101100: fc_kernel = 8'hea;
     14'b01000001101101: fc_kernel = 8'hec;
     14'b01000001101110: fc_kernel = 8'hed;
     14'b01000001101111: fc_kernel = 8'hf0;
     14'b01000001110000: fc_kernel = 8'hf0;
     14'b01000001110001: fc_kernel = 8'hfa;
     14'b01000001110010: fc_kernel = 8'hf7;
     14'b01000001110011: fc_kernel = 8'hf5;
     14'b01000001110100: fc_kernel = 8'h04;
     14'b01000001110101: fc_kernel = 8'h0b;
     14'b01000001110110: fc_kernel = 8'h04;
     14'b01000001110111: fc_kernel = 8'hf1;
     14'b01000001111000: fc_kernel = 8'hf2;
     14'b01000001111001: fc_kernel = 8'hfb;
     14'b01000001111010: fc_kernel = 8'h0e;
     14'b01000001111011: fc_kernel = 8'h0e;
     14'b01000001111100: fc_kernel = 8'h00;
     14'b01000001111101: fc_kernel = 8'hfd;
     14'b01000001111110: fc_kernel = 8'h00;
     14'b01000001111111: fc_kernel = 8'hfb;
     14'b01000010000000: fc_kernel = 8'hf5;
     14'b01000010000001: fc_kernel = 8'hf3;
     14'b01000010000010: fc_kernel = 8'he8;
     14'b01000010000011: fc_kernel = 8'hea;
     14'b01000010000100: fc_kernel = 8'he9;
     14'b01000010000101: fc_kernel = 8'heb;
     14'b01000010000110: fc_kernel = 8'hee;
     14'b01000010000111: fc_kernel = 8'hee;
     14'b01000010001000: fc_kernel = 8'hf1;
     14'b01000010001001: fc_kernel = 8'hf4;
     14'b01000010001010: fc_kernel = 8'hfb;
     14'b01000010001011: fc_kernel = 8'hf6;
     14'b01000010001100: fc_kernel = 8'hfd;
     14'b01000010001101: fc_kernel = 8'h05;
     14'b01000010001110: fc_kernel = 8'h05;
     14'b01000010001111: fc_kernel = 8'h01;
     14'b01000010010000: fc_kernel = 8'hf9;
     14'b01000010010001: fc_kernel = 8'hf7;
     14'b01000010010010: fc_kernel = 8'h07;
     14'b01000010010011: fc_kernel = 8'h05;
     14'b01000010010100: fc_kernel = 8'h00;
     14'b01000010010101: fc_kernel = 8'hfe;
     14'b01000010010110: fc_kernel = 8'hf8;
     14'b01000010010111: fc_kernel = 8'hf8;
     14'b01000010011000: fc_kernel = 8'hf8;
     14'b01000010011001: fc_kernel = 8'hf0;
     14'b01000010011010: fc_kernel = 8'hed;
     14'b01000010011011: fc_kernel = 8'hed;
     14'b01000010011100: fc_kernel = 8'hed;
     14'b01000010011101: fc_kernel = 8'heb;
     14'b01000010011110: fc_kernel = 8'hee;
     14'b01000010011111: fc_kernel = 8'hf0;
     14'b01000010100000: fc_kernel = 8'hf7;
     14'b01000010100001: fc_kernel = 8'hf7;
     14'b01000010100010: fc_kernel = 8'hfb;
     14'b01000010100011: fc_kernel = 8'hf4;
     14'b01000010100100: fc_kernel = 8'hfd;
     14'b01000010100101: fc_kernel = 8'hfb;
     14'b01000010100110: fc_kernel = 8'hfe;
     14'b01000010100111: fc_kernel = 8'hff;
     14'b01000010101000: fc_kernel = 8'hec;
     14'b01000010101001: fc_kernel = 8'hed;
     14'b01000010101010: fc_kernel = 8'hf8;
     14'b01000010101011: fc_kernel = 8'hf4;
     14'b01000010101100: fc_kernel = 8'hfd;
     14'b01000010101101: fc_kernel = 8'hfc;
     14'b01000010101110: fc_kernel = 8'hfe;
     14'b01000010101111: fc_kernel = 8'hf4;
     14'b01000010110000: fc_kernel = 8'hf9;
     14'b01000010110001: fc_kernel = 8'hf3;
     14'b01000010110010: fc_kernel = 8'hf7;
     14'b01000010110011: fc_kernel = 8'hf0;
     14'b01000010110100: fc_kernel = 8'hec;
     14'b01000010110101: fc_kernel = 8'hea;
     14'b01000010110110: fc_kernel = 8'hef;
     14'b01000010110111: fc_kernel = 8'hf4;
     14'b01000010111000: fc_kernel = 8'hf6;
     14'b01000010111001: fc_kernel = 8'h00;
     14'b01000010111010: fc_kernel = 8'hfe;
     14'b01000010111011: fc_kernel = 8'hfc;
     14'b01000010111100: fc_kernel = 8'hf8;
     14'b01000010111101: fc_kernel = 8'hf6;
     14'b01000010111110: fc_kernel = 8'hf1;
     14'b01000010111111: fc_kernel = 8'hf2;
     14'b01000011000000: fc_kernel = 8'he9;
     14'b01000011000001: fc_kernel = 8'hef;
     14'b01000011000010: fc_kernel = 8'hfa;
     14'b01000011000011: fc_kernel = 8'hf5;
     14'b01000011000100: fc_kernel = 8'hf5;
     14'b01000011000101: fc_kernel = 8'hf2;
     14'b01000011000110: fc_kernel = 8'hfe;
     14'b01000011000111: fc_kernel = 8'hfe;
     14'b01000011001000: fc_kernel = 8'hfa;
     14'b01000011001001: fc_kernel = 8'hf8;
     14'b01000011001010: fc_kernel = 8'hfc;
     14'b01000011001011: fc_kernel = 8'heb;
     14'b01000011001100: fc_kernel = 8'hdc;
     14'b01000011001101: fc_kernel = 8'he8;
     14'b01000011001110: fc_kernel = 8'hfe;
     14'b01000011001111: fc_kernel = 8'h00;
     14'b01000011010000: fc_kernel = 8'h00;
     14'b01000011010001: fc_kernel = 8'h00;
     14'b01000011010010: fc_kernel = 8'hf9;
     14'b01000011010011: fc_kernel = 8'hfe;
     14'b01000011010100: fc_kernel = 8'hf7;
     14'b01000011010101: fc_kernel = 8'hec;
     14'b01000011010110: fc_kernel = 8'he3;
     14'b01000011010111: fc_kernel = 8'hdb;
     14'b01000011011000: fc_kernel = 8'he9;
     14'b01000011011001: fc_kernel = 8'hf1;
     14'b01000011011010: fc_kernel = 8'hf6;
     14'b01000011011011: fc_kernel = 8'hf4;
     14'b01000011011100: fc_kernel = 8'hfc;
     14'b01000011011101: fc_kernel = 8'hf5;
     14'b01000011011110: fc_kernel = 8'h05;
     14'b01000011011111: fc_kernel = 8'h07;
     14'b01000011100000: fc_kernel = 8'h07;
     14'b01000011100001: fc_kernel = 8'h08;
     14'b01000011100010: fc_kernel = 8'h0a;
     14'b01000011100011: fc_kernel = 8'heb;
     14'b01000011100100: fc_kernel = 8'hde;
     14'b01000011100101: fc_kernel = 8'hf3;
     14'b01000011100110: fc_kernel = 8'h08;
     14'b01000011100111: fc_kernel = 8'h00;
     14'b01000011101000: fc_kernel = 8'h00;
     14'b01000011101001: fc_kernel = 8'hfd;
     14'b01000011101010: fc_kernel = 8'hfa;
     14'b01000011101011: fc_kernel = 8'hf9;
     14'b01000011101100: fc_kernel = 8'hf6;
     14'b01000011101101: fc_kernel = 8'heb;
     14'b01000011101110: fc_kernel = 8'hd7;
     14'b01000011101111: fc_kernel = 8'hd0;
     14'b01000011110000: fc_kernel = 8'hf0;
     14'b01000011110001: fc_kernel = 8'hee;
     14'b01000011110010: fc_kernel = 8'he9;
     14'b01000011110011: fc_kernel = 8'hf6;
     14'b01000011110100: fc_kernel = 8'h00;
     14'b01000011110101: fc_kernel = 8'h07;
     14'b01000011110110: fc_kernel = 8'h09;
     14'b01000011110111: fc_kernel = 8'h0f;
     14'b01000011111000: fc_kernel = 8'h10;
     14'b01000011111001: fc_kernel = 8'h17;
     14'b01000011111010: fc_kernel = 8'h13;
     14'b01000011111011: fc_kernel = 8'hfb;
     14'b01000011111100: fc_kernel = 8'he5;
     14'b01000011111101: fc_kernel = 8'hfd;
     14'b01000011111110: fc_kernel = 8'h0c;
     14'b01000011111111: fc_kernel = 8'h07;
     14'b01000100000000: fc_kernel = 8'h00;
     14'b01000100000001: fc_kernel = 8'hff;
     14'b01000100000010: fc_kernel = 8'h02;
     14'b01000100000011: fc_kernel = 8'hfe;
     14'b01000100000100: fc_kernel = 8'hfa;
     14'b01000100000101: fc_kernel = 8'hee;
     14'b01000100000110: fc_kernel = 8'he7;
     14'b01000100000111: fc_kernel = 8'hdf;
     14'b01000100001000: fc_kernel = 8'hed;
     14'b01000100001001: fc_kernel = 8'hf3;
     14'b01000100001010: fc_kernel = 8'hfb;
     14'b01000100001011: fc_kernel = 8'h00;
     14'b01000100001100: fc_kernel = 8'h0e;
     14'b01000100001101: fc_kernel = 8'h0d;
     14'b01000100001110: fc_kernel = 8'h10;
     14'b01000100001111: fc_kernel = 8'h0c;
     14'b01000100010000: fc_kernel = 8'h0f;
     14'b01000100010001: fc_kernel = 8'h1a;
     14'b01000100010010: fc_kernel = 8'h11;
     14'b01000100010011: fc_kernel = 8'hf9;
     14'b01000100010100: fc_kernel = 8'hf4;
     14'b01000100010101: fc_kernel = 8'h08;
     14'b01000100010110: fc_kernel = 8'h0e;
     14'b01000100010111: fc_kernel = 8'h0e;
     14'b01000100011000: fc_kernel = 8'h02;
     14'b01000100011001: fc_kernel = 8'h07;
     14'b01000100011010: fc_kernel = 8'h0e;
     14'b01000100011011: fc_kernel = 8'h0f;
     14'b01000100011100: fc_kernel = 8'h07;
     14'b01000100011101: fc_kernel = 8'h00;
     14'b01000100011110: fc_kernel = 8'hf9;
     14'b01000100011111: fc_kernel = 8'hf5;
     14'b01000100100000: fc_kernel = 8'hea;
     14'b01000100100001: fc_kernel = 8'h07;
     14'b01000100100010: fc_kernel = 8'h09;
     14'b01000100100011: fc_kernel = 8'h12;
     14'b01000100100100: fc_kernel = 8'h0f;
     14'b01000100100101: fc_kernel = 8'h0c;
     14'b01000100100110: fc_kernel = 8'h12;
     14'b01000100100111: fc_kernel = 8'h0a;
     14'b01000100101000: fc_kernel = 8'h12;
     14'b01000100101001: fc_kernel = 8'h14;
     14'b01000100101010: fc_kernel = 8'h0f;
     14'b01000100101011: fc_kernel = 8'hf7;
     14'b01000100101100: fc_kernel = 8'hfa;
     14'b01000100101101: fc_kernel = 8'h0c;
     14'b01000100101110: fc_kernel = 8'h0f;
     14'b01000100101111: fc_kernel = 8'h11;
     14'b01000100110000: fc_kernel = 8'h0f;
     14'b01000100110001: fc_kernel = 8'h04;
     14'b01000100110010: fc_kernel = 8'h06;
     14'b01000100110011: fc_kernel = 8'h0b;
     14'b01000100110100: fc_kernel = 8'h06;
     14'b01000100110101: fc_kernel = 8'hf6;
     14'b01000100110110: fc_kernel = 8'heb;
     14'b01000100110111: fc_kernel = 8'he9;
     14'b01000100111000: fc_kernel = 8'hf0;
     14'b01000100111001: fc_kernel = 8'h0a;
     14'b01000100111010: fc_kernel = 8'h0f;
     14'b01000100111011: fc_kernel = 8'h0c;
     14'b01000100111100: fc_kernel = 8'h0c;
     14'b01000100111101: fc_kernel = 8'h0c;
     14'b01000100111110: fc_kernel = 8'h0c;
     14'b01000100111111: fc_kernel = 8'h09;
     14'b01000101000000: fc_kernel = 8'h10;
     14'b01000101000001: fc_kernel = 8'h14;
     14'b01000101000010: fc_kernel = 8'h0d;
     14'b01000101000011: fc_kernel = 8'hfd;
     14'b01000101000100: fc_kernel = 8'hff;
     14'b01000101000101: fc_kernel = 8'h0c;
     14'b01000101000110: fc_kernel = 8'h15;
     14'b01000101000111: fc_kernel = 8'h10;
     14'b01000101001000: fc_kernel = 8'h0e;
     14'b01000101001001: fc_kernel = 8'h07;
     14'b01000101001010: fc_kernel = 8'h01;
     14'b01000101001011: fc_kernel = 8'h01;
     14'b01000101001100: fc_kernel = 8'h01;
     14'b01000101001101: fc_kernel = 8'hf7;
     14'b01000101001110: fc_kernel = 8'he3;
     14'b01000101001111: fc_kernel = 8'hdd;
     14'b01000101010000: fc_kernel = 8'hfa;
     14'b01000101010001: fc_kernel = 8'h00;
     14'b01000101010010: fc_kernel = 8'hf9;
     14'b01000101010011: fc_kernel = 8'hfb;
     14'b01000101010100: fc_kernel = 8'h01;
     14'b01000101010101: fc_kernel = 8'h0d;
     14'b01000101010110: fc_kernel = 8'h0c;
     14'b01000101010111: fc_kernel = 8'h09;
     14'b01000101011000: fc_kernel = 8'h08;
     14'b01000101011001: fc_kernel = 8'h01;
     14'b01000101011010: fc_kernel = 8'hfc;
     14'b01000101011011: fc_kernel = 8'hfb;
     14'b01000101011100: fc_kernel = 8'h02;
     14'b01000101011101: fc_kernel = 8'h16;
     14'b01000101011110: fc_kernel = 8'h1d;
     14'b01000101011111: fc_kernel = 8'h0d;
     14'b01000101100000: fc_kernel = 8'h0b;
     14'b01000101100001: fc_kernel = 8'h05;
     14'b01000101100010: fc_kernel = 8'h04;
     14'b01000101100011: fc_kernel = 8'h00;
     14'b01000101100100: fc_kernel = 8'h02;
     14'b01000101100101: fc_kernel = 8'hf8;
     14'b01000101100110: fc_kernel = 8'he5;
     14'b01000101100111: fc_kernel = 8'hd7;
     14'b01000101101000: fc_kernel = 8'hf6;
     14'b01000101101001: fc_kernel = 8'hed;
     14'b01000101101010: fc_kernel = 8'hed;
     14'b01000101101011: fc_kernel = 8'hf1;
     14'b01000101101100: fc_kernel = 8'hfd;
     14'b01000101101101: fc_kernel = 8'h0a;
     14'b01000101101110: fc_kernel = 8'h12;
     14'b01000101101111: fc_kernel = 8'h09;
     14'b01000101110000: fc_kernel = 8'h00;
     14'b01000101110001: fc_kernel = 8'h01;
     14'b01000101110010: fc_kernel = 8'h01;
     14'b01000101110011: fc_kernel = 8'h05;
     14'b01000101110100: fc_kernel = 8'h0f;
     14'b01000101110101: fc_kernel = 8'h18;
     14'b01000101110110: fc_kernel = 8'h11;
     14'b01000101110111: fc_kernel = 8'h0b;
     14'b01000101111000: fc_kernel = 8'h05;
     14'b01000101111001: fc_kernel = 8'h00;
     14'b01000101111010: fc_kernel = 8'h05;
     14'b01000101111011: fc_kernel = 8'h09;
     14'b01000101111100: fc_kernel = 8'h01;
     14'b01000101111101: fc_kernel = 8'hf9;
     14'b01000101111110: fc_kernel = 8'he7;
     14'b01000101111111: fc_kernel = 8'hda;
     14'b01000110000000: fc_kernel = 8'hf3;
     14'b01000110000001: fc_kernel = 8'heb;
     14'b01000110000010: fc_kernel = 8'hf0;
     14'b01000110000011: fc_kernel = 8'hfa;
     14'b01000110000100: fc_kernel = 8'h04;
     14'b01000110000101: fc_kernel = 8'h03;
     14'b01000110000110: fc_kernel = 8'h08;
     14'b01000110000111: fc_kernel = 8'h06;
     14'b01000110001000: fc_kernel = 8'hfe;
     14'b01000110001001: fc_kernel = 8'hfb;
     14'b01000110001010: fc_kernel = 8'h00;
     14'b01000110001011: fc_kernel = 8'h09;
     14'b01000110001100: fc_kernel = 8'h12;
     14'b01000110001101: fc_kernel = 8'h0f;
     14'b01000110001110: fc_kernel = 8'h0d;
     14'b01000110001111: fc_kernel = 8'h05;
     14'b01000110010000: fc_kernel = 8'hfe;
     14'b01000110010001: fc_kernel = 8'h00;
     14'b01000110010010: fc_kernel = 8'hff;
     14'b01000110010011: fc_kernel = 8'h00;
     14'b01000110010100: fc_kernel = 8'hfb;
     14'b01000110010101: fc_kernel = 8'hf0;
     14'b01000110010110: fc_kernel = 8'hec;
     14'b01000110010111: fc_kernel = 8'hd7;
     14'b01000110011000: fc_kernel = 8'hf9;
     14'b01000110011001: fc_kernel = 8'hfb;
     14'b01000110011010: fc_kernel = 8'hfd;
     14'b01000110011011: fc_kernel = 8'hf9;
     14'b01000110011100: fc_kernel = 8'hfe;
     14'b01000110011101: fc_kernel = 8'h01;
     14'b01000110011110: fc_kernel = 8'hfa;
     14'b01000110011111: fc_kernel = 8'hf3;
     14'b01000110100000: fc_kernel = 8'hec;
     14'b01000110100001: fc_kernel = 8'hed;
     14'b01000110100010: fc_kernel = 8'hf7;
     14'b01000110100011: fc_kernel = 8'h02;
     14'b01000110100100: fc_kernel = 8'h0b;
     14'b01000110100101: fc_kernel = 8'h0e;
     14'b01000110100110: fc_kernel = 8'h05;
     14'b01000110100111: fc_kernel = 8'h03;
     14'b01000110101000: fc_kernel = 8'hfa;
     14'b01000110101001: fc_kernel = 8'hf8;
     14'b01000110101010: fc_kernel = 8'hfb;
     14'b01000110101011: fc_kernel = 8'hfa;
     14'b01000110101100: fc_kernel = 8'hee;
     14'b01000110101101: fc_kernel = 8'he4;
     14'b01000110101110: fc_kernel = 8'he1;
     14'b01000110101111: fc_kernel = 8'hd1;
     14'b01000110110000: fc_kernel = 8'h00;
     14'b01000110110001: fc_kernel = 8'h03;
     14'b01000110110010: fc_kernel = 8'hf8;
     14'b01000110110011: fc_kernel = 8'h00;
     14'b01000110110100: fc_kernel = 8'hfe;
     14'b01000110110101: fc_kernel = 8'hf9;
     14'b01000110110110: fc_kernel = 8'hf8;
     14'b01000110110111: fc_kernel = 8'hf2;
     14'b01000110111000: fc_kernel = 8'hf4;
     14'b01000110111001: fc_kernel = 8'hf1;
     14'b01000110111010: fc_kernel = 8'hf6;
     14'b01000110111011: fc_kernel = 8'hfa;
     14'b01000110111100: fc_kernel = 8'h02;
     14'b01000110111101: fc_kernel = 8'h0e;
     14'b01000110111110: fc_kernel = 8'h04;
     14'b01000110111111: fc_kernel = 8'hfe;
     14'b01000111000000: fc_kernel = 8'h00;
     14'b01000111000001: fc_kernel = 8'hfc;
     14'b01000111000010: fc_kernel = 8'hfa;
     14'b01000111000011: fc_kernel = 8'hf5;
     14'b01000111000100: fc_kernel = 8'hed;
     14'b01000111000101: fc_kernel = 8'he0;
     14'b01000111000110: fc_kernel = 8'hdf;
     14'b01000111000111: fc_kernel = 8'hd7;
     14'b01000111001000: fc_kernel = 8'hfd;
     14'b01000111001001: fc_kernel = 8'hf8;
     14'b01000111001010: fc_kernel = 8'hfb;
     14'b01000111001011: fc_kernel = 8'hf4;
     14'b01000111001100: fc_kernel = 8'hf0;
     14'b01000111001101: fc_kernel = 8'hed;
     14'b01000111001110: fc_kernel = 8'heb;
     14'b01000111001111: fc_kernel = 8'hf0;
     14'b01000111010000: fc_kernel = 8'hf6;
     14'b01000111010001: fc_kernel = 8'hf2;
     14'b01000111010010: fc_kernel = 8'hf5;
     14'b01000111010011: fc_kernel = 8'hf9;
     14'b01000111010100: fc_kernel = 8'h00;
     14'b01000111010101: fc_kernel = 8'hfe;
     14'b01000111010110: fc_kernel = 8'hfe;
     14'b01000111010111: fc_kernel = 8'hfe;
     14'b01000111011000: fc_kernel = 8'hfb;
     14'b01000111011001: fc_kernel = 8'hfc;
     14'b01000111011010: fc_kernel = 8'h00;
     14'b01000111011011: fc_kernel = 8'hfb;
     14'b01000111011100: fc_kernel = 8'hfe;
     14'b01000111011101: fc_kernel = 8'hfa;
     14'b01000111011110: fc_kernel = 8'hed;
     14'b01000111011111: fc_kernel = 8'he2;
     14'b01000111100000: fc_kernel = 8'hef;
     14'b01000111100001: fc_kernel = 8'hed;
     14'b01000111100010: fc_kernel = 8'he5;
     14'b01000111100011: fc_kernel = 8'heb;
     14'b01000111100100: fc_kernel = 8'he9;
     14'b01000111100101: fc_kernel = 8'hf1;
     14'b01000111100110: fc_kernel = 8'hf8;
     14'b01000111100111: fc_kernel = 8'hf6;
     14'b01000111101000: fc_kernel = 8'hf7;
     14'b01000111101001: fc_kernel = 8'hfe;
     14'b01000111101010: fc_kernel = 8'hfd;
     14'b01000111101011: fc_kernel = 8'hfb;
     14'b01000111101100: fc_kernel = 8'h01;
     14'b01000111101101: fc_kernel = 8'h01;
     14'b01000111101110: fc_kernel = 8'h01;
     14'b01000111101111: fc_kernel = 8'h01;
     14'b01000111110000: fc_kernel = 8'h00;
     14'b01000111110001: fc_kernel = 8'hfe;
     14'b01000111110010: fc_kernel = 8'h05;
     14'b01000111110011: fc_kernel = 8'h00;
     14'b01000111110100: fc_kernel = 8'hfb;
     14'b01000111110101: fc_kernel = 8'hff;
     14'b01000111110110: fc_kernel = 8'hf3;
     14'b01000111110111: fc_kernel = 8'hed;
     14'b01000111111000: fc_kernel = 8'heb;
     14'b01000111111001: fc_kernel = 8'hdf;
     14'b01000111111010: fc_kernel = 8'hd9;
     14'b01000111111011: fc_kernel = 8'hea;
     14'b01000111111100: fc_kernel = 8'hff;
     14'b01000111111101: fc_kernel = 8'h05;
     14'b01000111111110: fc_kernel = 8'h07;
     14'b01000111111111: fc_kernel = 8'hfe;
     14'b01001000000000: fc_kernel = 8'h04;
     14'b01001000000001: fc_kernel = 8'h03;
     14'b01001000000010: fc_kernel = 8'h01;
     14'b01001000000011: fc_kernel = 8'h03;
     14'b01001000000100: fc_kernel = 8'h05;
     14'b01001000000101: fc_kernel = 8'h02;
     14'b01001000000110: fc_kernel = 8'h06;
     14'b01001000000111: fc_kernel = 8'h05;
     14'b01001000001000: fc_kernel = 8'h0e;
     14'b01001000001001: fc_kernel = 8'h09;
     14'b01001000001010: fc_kernel = 8'h0a;
     14'b01001000001011: fc_kernel = 8'h0a;
     14'b01001000001100: fc_kernel = 8'h05;
     14'b01001000001101: fc_kernel = 8'hfa;
     14'b01001000001110: fc_kernel = 8'hf1;
     14'b01001000001111: fc_kernel = 8'hf6;
     14'b01001000010000: fc_kernel = 8'he4;
     14'b01001000010001: fc_kernel = 8'he3;
     14'b01001000010010: fc_kernel = 8'hd5;
     14'b01001000010011: fc_kernel = 8'hf0;
     14'b01001000010100: fc_kernel = 8'h00;
     14'b01001000010101: fc_kernel = 8'h02;
     14'b01001000010110: fc_kernel = 8'h01;
     14'b01001000010111: fc_kernel = 8'h02;
     14'b01001000011000: fc_kernel = 8'h08;
     14'b01001000011001: fc_kernel = 8'h03;
     14'b01001000011010: fc_kernel = 8'h04;
     14'b01001000011011: fc_kernel = 8'h04;
     14'b01001000011100: fc_kernel = 8'h05;
     14'b01001000011101: fc_kernel = 8'h08;
     14'b01001000011110: fc_kernel = 8'h07;
     14'b01001000011111: fc_kernel = 8'h00;
     14'b01001000100000: fc_kernel = 8'h02;
     14'b01001000100001: fc_kernel = 8'h05;
     14'b01001000100010: fc_kernel = 8'h09;
     14'b01001000100011: fc_kernel = 8'h05;
     14'b01001000100100: fc_kernel = 8'h00;
     14'b01001000100101: fc_kernel = 8'hfe;
     14'b01001000100110: fc_kernel = 8'hf6;
     14'b01001000100111: fc_kernel = 8'hf6;
     14'b01001000101000: fc_kernel = 8'he7;
     14'b01001000101001: fc_kernel = 8'hf2;
     14'b01001000101010: fc_kernel = 8'hf4;
     14'b01001000101011: fc_kernel = 8'hf8;
     14'b01001000101100: fc_kernel = 8'hf8;
     14'b01001000101101: fc_kernel = 8'hf1;
     14'b01001000101110: fc_kernel = 8'he7;
     14'b01001000101111: fc_kernel = 8'hea;
     14'b01001000110000: fc_kernel = 8'hf6;
     14'b01001000110001: fc_kernel = 8'hea;
     14'b01001000110010: fc_kernel = 8'he5;
     14'b01001000110011: fc_kernel = 8'he3;
     14'b01001000110100: fc_kernel = 8'heb;
     14'b01001000110101: fc_kernel = 8'he9;
     14'b01001000110110: fc_kernel = 8'he8;
     14'b01001000110111: fc_kernel = 8'he4;
     14'b01001000111000: fc_kernel = 8'he2;
     14'b01001000111001: fc_kernel = 8'he9;
     14'b01001000111010: fc_kernel = 8'hec;
     14'b01001000111011: fc_kernel = 8'hf6;
     14'b01001000111100: fc_kernel = 8'hfc;
     14'b01001000111101: fc_kernel = 8'hfb;
     14'b01001000111110: fc_kernel = 8'hf4;
     14'b01001000111111: fc_kernel = 8'hf8;
     14'b01010000000000: fc_kernel = 8'he4;
     14'b01010000000001: fc_kernel = 8'hf4;
     14'b01010000000010: fc_kernel = 8'h08;
     14'b01010000000011: fc_kernel = 8'h07;
     14'b01010000000100: fc_kernel = 8'he9;
     14'b01010000000101: fc_kernel = 8'h16;
     14'b01010000000110: fc_kernel = 8'hfa;
     14'b01010000000111: fc_kernel = 8'hfd;
     14'b01010000001000: fc_kernel = 8'hdc;
     14'b01010000001001: fc_kernel = 8'hd9;
     14'b01010000001010: fc_kernel = 8'hd9;
     14'b01010000001011: fc_kernel = 8'hdb;
     14'b01010000001100: fc_kernel = 8'he0;
     14'b01010000001101: fc_kernel = 8'hed;
     14'b01010000001110: fc_kernel = 8'hfd;
     14'b01010000001111: fc_kernel = 8'h07;
     14'b01010000010000: fc_kernel = 8'h10;
     14'b01010000010001: fc_kernel = 8'h10;
     14'b01010000010010: fc_kernel = 8'h08;
     14'b01010000010011: fc_kernel = 8'h03;
     14'b01010000010100: fc_kernel = 8'hf8;
     14'b01010000010101: fc_kernel = 8'hf2;
     14'b01010000010110: fc_kernel = 8'hf5;
     14'b01010000010111: fc_kernel = 8'h01;
     14'b01010000011000: fc_kernel = 8'he0;
     14'b01010000011001: fc_kernel = 8'h08;
     14'b01010000011010: fc_kernel = 8'hfa;
     14'b01010000011011: fc_kernel = 8'h03;
     14'b01010000011100: fc_kernel = 8'h05;
     14'b01010000011101: fc_kernel = 8'h00;
     14'b01010000011110: fc_kernel = 8'hfb;
     14'b01010000011111: fc_kernel = 8'hfe;
     14'b01010000100000: fc_kernel = 8'hfd;
     14'b01010000100001: fc_kernel = 8'hf4;
     14'b01010000100010: fc_kernel = 8'hf8;
     14'b01010000100011: fc_kernel = 8'hfa;
     14'b01010000100100: fc_kernel = 8'hff;
     14'b01010000100101: fc_kernel = 8'h07;
     14'b01010000100110: fc_kernel = 8'h04;
     14'b01010000100111: fc_kernel = 8'h05;
     14'b01010000101000: fc_kernel = 8'h11;
     14'b01010000101001: fc_kernel = 8'h09;
     14'b01010000101010: fc_kernel = 8'h13;
     14'b01010000101011: fc_kernel = 8'h1a;
     14'b01010000101100: fc_kernel = 8'h13;
     14'b01010000101101: fc_kernel = 8'h02;
     14'b01010000101110: fc_kernel = 8'h01;
     14'b01010000101111: fc_kernel = 8'h0b;
     14'b01010000110000: fc_kernel = 8'h01;
     14'b01010000110001: fc_kernel = 8'h07;
     14'b01010000110010: fc_kernel = 8'hd8;
     14'b01010000110011: fc_kernel = 8'he8;
     14'b01010000110100: fc_kernel = 8'hf2;
     14'b01010000110101: fc_kernel = 8'hf5;
     14'b01010000110110: fc_kernel = 8'hf5;
     14'b01010000110111: fc_kernel = 8'hf9;
     14'b01010000111000: fc_kernel = 8'h03;
     14'b01010000111001: fc_kernel = 8'h08;
     14'b01010000111010: fc_kernel = 8'h01;
     14'b01010000111011: fc_kernel = 8'h00;
     14'b01010000111100: fc_kernel = 8'h00;
     14'b01010000111101: fc_kernel = 8'h0c;
     14'b01010000111110: fc_kernel = 8'h0a;
     14'b01010000111111: fc_kernel = 8'h0c;
     14'b01010001000000: fc_kernel = 8'h0a;
     14'b01010001000001: fc_kernel = 8'h08;
     14'b01010001000010: fc_kernel = 8'h03;
     14'b01010001000011: fc_kernel = 8'h0e;
     14'b01010001000100: fc_kernel = 8'h0f;
     14'b01010001000101: fc_kernel = 8'h0d;
     14'b01010001000110: fc_kernel = 8'h11;
     14'b01010001000111: fc_kernel = 8'h1e;
     14'b01010001001000: fc_kernel = 8'he0;
     14'b01010001001001: fc_kernel = 8'hef;
     14'b01010001001010: fc_kernel = 8'hea;
     14'b01010001001011: fc_kernel = 8'hed;
     14'b01010001001100: fc_kernel = 8'hf4;
     14'b01010001001101: fc_kernel = 8'hf8;
     14'b01010001001110: fc_kernel = 8'hfb;
     14'b01010001001111: fc_kernel = 8'hfd;
     14'b01010001010000: fc_kernel = 8'h05;
     14'b01010001010001: fc_kernel = 8'h03;
     14'b01010001010010: fc_kernel = 8'h00;
     14'b01010001010011: fc_kernel = 8'hfc;
     14'b01010001010100: fc_kernel = 8'hff;
     14'b01010001010101: fc_kernel = 8'h04;
     14'b01010001010110: fc_kernel = 8'h02;
     14'b01010001010111: fc_kernel = 8'h0a;
     14'b01010001011000: fc_kernel = 8'h0d;
     14'b01010001011001: fc_kernel = 8'h06;
     14'b01010001011010: fc_kernel = 8'h09;
     14'b01010001011011: fc_kernel = 8'h08;
     14'b01010001011100: fc_kernel = 8'h0b;
     14'b01010001011101: fc_kernel = 8'h14;
     14'b01010001011110: fc_kernel = 8'h14;
     14'b01010001011111: fc_kernel = 8'h24;
     14'b01010001100000: fc_kernel = 8'hd2;
     14'b01010001100001: fc_kernel = 8'he3;
     14'b01010001100010: fc_kernel = 8'hed;
     14'b01010001100011: fc_kernel = 8'hf9;
     14'b01010001100100: fc_kernel = 8'h05;
     14'b01010001100101: fc_kernel = 8'h01;
     14'b01010001100110: fc_kernel = 8'hfe;
     14'b01010001100111: fc_kernel = 8'h02;
     14'b01010001101000: fc_kernel = 8'h00;
     14'b01010001101001: fc_kernel = 8'h00;
     14'b01010001101010: fc_kernel = 8'h00;
     14'b01010001101011: fc_kernel = 8'h04;
     14'b01010001101100: fc_kernel = 8'h01;
     14'b01010001101101: fc_kernel = 8'h02;
     14'b01010001101110: fc_kernel = 8'h04;
     14'b01010001101111: fc_kernel = 8'h07;
     14'b01010001110000: fc_kernel = 8'h06;
     14'b01010001110001: fc_kernel = 8'h0b;
     14'b01010001110010: fc_kernel = 8'h06;
     14'b01010001110011: fc_kernel = 8'h08;
     14'b01010001110100: fc_kernel = 8'h04;
     14'b01010001110101: fc_kernel = 8'h0d;
     14'b01010001110110: fc_kernel = 8'h17;
     14'b01010001110111: fc_kernel = 8'h30;
     14'b01010001111000: fc_kernel = 8'he6;
     14'b01010001111001: fc_kernel = 8'hd0;
     14'b01010001111010: fc_kernel = 8'hdf;
     14'b01010001111011: fc_kernel = 8'hfa;
     14'b01010001111100: fc_kernel = 8'h02;
     14'b01010001111101: fc_kernel = 8'hfd;
     14'b01010001111110: fc_kernel = 8'h07;
     14'b01010001111111: fc_kernel = 8'h03;
     14'b01010010000000: fc_kernel = 8'h00;
     14'b01010010000001: fc_kernel = 8'h07;
     14'b01010010000010: fc_kernel = 8'h00;
     14'b01010010000011: fc_kernel = 8'h00;
     14'b01010010000100: fc_kernel = 8'h04;
     14'b01010010000101: fc_kernel = 8'h02;
     14'b01010010000110: fc_kernel = 8'h09;
     14'b01010010000111: fc_kernel = 8'h07;
     14'b01010010001000: fc_kernel = 8'h05;
     14'b01010010001001: fc_kernel = 8'h0c;
     14'b01010010001010: fc_kernel = 8'h04;
     14'b01010010001011: fc_kernel = 8'h06;
     14'b01010010001100: fc_kernel = 8'h05;
     14'b01010010001101: fc_kernel = 8'h0e;
     14'b01010010001110: fc_kernel = 8'h1e;
     14'b01010010001111: fc_kernel = 8'h2d;
     14'b01010010010000: fc_kernel = 8'he3;
     14'b01010010010001: fc_kernel = 8'hca;
     14'b01010010010010: fc_kernel = 8'he1;
     14'b01010010010011: fc_kernel = 8'hf2;
     14'b01010010010100: fc_kernel = 8'hfc;
     14'b01010010010101: fc_kernel = 8'hfb;
     14'b01010010010110: fc_kernel = 8'h00;
     14'b01010010010111: fc_kernel = 8'h00;
     14'b01010010011000: fc_kernel = 8'h04;
     14'b01010010011001: fc_kernel = 8'h06;
     14'b01010010011010: fc_kernel = 8'h01;
     14'b01010010011011: fc_kernel = 8'hfd;
     14'b01010010011100: fc_kernel = 8'hfe;
     14'b01010010011101: fc_kernel = 8'hfa;
     14'b01010010011110: fc_kernel = 8'h00;
     14'b01010010011111: fc_kernel = 8'h01;
     14'b01010010100000: fc_kernel = 8'h03;
     14'b01010010100001: fc_kernel = 8'h07;
     14'b01010010100010: fc_kernel = 8'h09;
     14'b01010010100011: fc_kernel = 8'h09;
     14'b01010010100100: fc_kernel = 8'h0e;
     14'b01010010100101: fc_kernel = 8'h11;
     14'b01010010100110: fc_kernel = 8'h25;
     14'b01010010100111: fc_kernel = 8'h2f;
     14'b01010010101000: fc_kernel = 8'hd8;
     14'b01010010101001: fc_kernel = 8'he0;
     14'b01010010101010: fc_kernel = 8'he9;
     14'b01010010101011: fc_kernel = 8'hf6;
     14'b01010010101100: fc_kernel = 8'hfe;
     14'b01010010101101: fc_kernel = 8'hfe;
     14'b01010010101110: fc_kernel = 8'h00;
     14'b01010010101111: fc_kernel = 8'h03;
     14'b01010010110000: fc_kernel = 8'h0a;
     14'b01010010110001: fc_kernel = 8'h0d;
     14'b01010010110010: fc_kernel = 8'h08;
     14'b01010010110011: fc_kernel = 8'h05;
     14'b01010010110100: fc_kernel = 8'hf6;
     14'b01010010110101: fc_kernel = 8'hf7;
     14'b01010010110110: fc_kernel = 8'hf5;
     14'b01010010110111: fc_kernel = 8'hf7;
     14'b01010010111000: fc_kernel = 8'hfe;
     14'b01010010111001: fc_kernel = 8'hfe;
     14'b01010010111010: fc_kernel = 8'h06;
     14'b01010010111011: fc_kernel = 8'h0e;
     14'b01010010111100: fc_kernel = 8'h0c;
     14'b01010010111101: fc_kernel = 8'h15;
     14'b01010010111110: fc_kernel = 8'h2c;
     14'b01010010111111: fc_kernel = 8'h3d;
     14'b01010011000000: fc_kernel = 8'hc0;
     14'b01010011000001: fc_kernel = 8'hea;
     14'b01010011000010: fc_kernel = 8'hef;
     14'b01010011000011: fc_kernel = 8'hf7;
     14'b01010011000100: fc_kernel = 8'hf9;
     14'b01010011000101: fc_kernel = 8'hff;
     14'b01010011000110: fc_kernel = 8'h07;
     14'b01010011000111: fc_kernel = 8'h0c;
     14'b01010011001000: fc_kernel = 8'h0b;
     14'b01010011001001: fc_kernel = 8'h0e;
     14'b01010011001010: fc_kernel = 8'h10;
     14'b01010011001011: fc_kernel = 8'h0a;
     14'b01010011001100: fc_kernel = 8'h00;
     14'b01010011001101: fc_kernel = 8'hf9;
     14'b01010011001110: fc_kernel = 8'hf6;
     14'b01010011001111: fc_kernel = 8'hf6;
     14'b01010011010000: fc_kernel = 8'hf4;
     14'b01010011010001: fc_kernel = 8'hf6;
     14'b01010011010010: fc_kernel = 8'hfc;
     14'b01010011010011: fc_kernel = 8'h04;
     14'b01010011010100: fc_kernel = 8'h06;
     14'b01010011010101: fc_kernel = 8'h24;
     14'b01010011010110: fc_kernel = 8'h3d;
     14'b01010011010111: fc_kernel = 8'h5a;
     14'b01010011011000: fc_kernel = 8'hc5;
     14'b01010011011001: fc_kernel = 8'hde;
     14'b01010011011010: fc_kernel = 8'hf4;
     14'b01010011011011: fc_kernel = 8'hf9;
     14'b01010011011100: fc_kernel = 8'h00;
     14'b01010011011101: fc_kernel = 8'h0b;
     14'b01010011011110: fc_kernel = 8'h0b;
     14'b01010011011111: fc_kernel = 8'h0d;
     14'b01010011100000: fc_kernel = 8'h0c;
     14'b01010011100001: fc_kernel = 8'h05;
     14'b01010011100010: fc_kernel = 8'h0c;
     14'b01010011100011: fc_kernel = 8'h0b;
     14'b01010011100100: fc_kernel = 8'h03;
     14'b01010011100101: fc_kernel = 8'hfc;
     14'b01010011100110: fc_kernel = 8'hfa;
     14'b01010011100111: fc_kernel = 8'hf7;
     14'b01010011101000: fc_kernel = 8'hf3;
     14'b01010011101001: fc_kernel = 8'hed;
     14'b01010011101010: fc_kernel = 8'heb;
     14'b01010011101011: fc_kernel = 8'he5;
     14'b01010011101100: fc_kernel = 8'hed;
     14'b01010011101101: fc_kernel = 8'h0b;
     14'b01010011101110: fc_kernel = 8'h34;
     14'b01010011101111: fc_kernel = 8'h5c;
     14'b01010011110000: fc_kernel = 8'hd4;
     14'b01010011110001: fc_kernel = 8'he3;
     14'b01010011110010: fc_kernel = 8'hf7;
     14'b01010011110011: fc_kernel = 8'h00;
     14'b01010011110100: fc_kernel = 8'h03;
     14'b01010011110101: fc_kernel = 8'h07;
     14'b01010011110110: fc_kernel = 8'h03;
     14'b01010011110111: fc_kernel = 8'h00;
     14'b01010011111000: fc_kernel = 8'h05;
     14'b01010011111001: fc_kernel = 8'h0c;
     14'b01010011111010: fc_kernel = 8'h0b;
     14'b01010011111011: fc_kernel = 8'h10;
     14'b01010011111100: fc_kernel = 8'hfe;
     14'b01010011111101: fc_kernel = 8'hf6;
     14'b01010011111110: fc_kernel = 8'hef;
     14'b01010011111111: fc_kernel = 8'hf7;
     14'b01010100000000: fc_kernel = 8'hf4;
     14'b01010100000001: fc_kernel = 8'hf8;
     14'b01010100000010: fc_kernel = 8'heb;
     14'b01010100000011: fc_kernel = 8'hdc;
     14'b01010100000100: fc_kernel = 8'hd3;
     14'b01010100000101: fc_kernel = 8'hd5;
     14'b01010100000110: fc_kernel = 8'hfb;
     14'b01010100000111: fc_kernel = 8'h24;
     14'b01010100001000: fc_kernel = 8'he2;
     14'b01010100001001: fc_kernel = 8'hfa;
     14'b01010100001010: fc_kernel = 8'h01;
     14'b01010100001011: fc_kernel = 8'h06;
     14'b01010100001100: fc_kernel = 8'h05;
     14'b01010100001101: fc_kernel = 8'h00;
     14'b01010100001110: fc_kernel = 8'hff;
     14'b01010100001111: fc_kernel = 8'hff;
     14'b01010100010000: fc_kernel = 8'h0b;
     14'b01010100010001: fc_kernel = 8'h0c;
     14'b01010100010010: fc_kernel = 8'h10;
     14'b01010100010011: fc_kernel = 8'h0b;
     14'b01010100010100: fc_kernel = 8'hff;
     14'b01010100010101: fc_kernel = 8'hf6;
     14'b01010100010110: fc_kernel = 8'hee;
     14'b01010100010111: fc_kernel = 8'hf4;
     14'b01010100011000: fc_kernel = 8'hf3;
     14'b01010100011001: fc_kernel = 8'hf8;
     14'b01010100011010: fc_kernel = 8'hf9;
     14'b01010100011011: fc_kernel = 8'hf2;
     14'b01010100011100: fc_kernel = 8'hdf;
     14'b01010100011101: fc_kernel = 8'hc9;
     14'b01010100011110: fc_kernel = 8'hbd;
     14'b01010100011111: fc_kernel = 8'hd8;
     14'b01010100100000: fc_kernel = 8'hef;
     14'b01010100100001: fc_kernel = 8'h05;
     14'b01010100100010: fc_kernel = 8'h04;
     14'b01010100100011: fc_kernel = 8'h03;
     14'b01010100100100: fc_kernel = 8'h00;
     14'b01010100100101: fc_kernel = 8'h04;
     14'b01010100100110: fc_kernel = 8'h00;
     14'b01010100100111: fc_kernel = 8'h08;
     14'b01010100101000: fc_kernel = 8'h09;
     14'b01010100101001: fc_kernel = 8'h0a;
     14'b01010100101010: fc_kernel = 8'h0b;
     14'b01010100101011: fc_kernel = 8'h00;
     14'b01010100101100: fc_kernel = 8'hfa;
     14'b01010100101101: fc_kernel = 8'hf3;
     14'b01010100101110: fc_kernel = 8'hf4;
     14'b01010100101111: fc_kernel = 8'hf1;
     14'b01010100110000: fc_kernel = 8'hfa;
     14'b01010100110001: fc_kernel = 8'hf6;
     14'b01010100110010: fc_kernel = 8'hf8;
     14'b01010100110011: fc_kernel = 8'hf4;
     14'b01010100110100: fc_kernel = 8'hf6;
     14'b01010100110101: fc_kernel = 8'hf1;
     14'b01010100110110: fc_kernel = 8'hdd;
     14'b01010100110111: fc_kernel = 8'hd2;
     14'b01010100111000: fc_kernel = 8'hfc;
     14'b01010100111001: fc_kernel = 8'h09;
     14'b01010100111010: fc_kernel = 8'h00;
     14'b01010100111011: fc_kernel = 8'hfa;
     14'b01010100111100: fc_kernel = 8'hf2;
     14'b01010100111101: fc_kernel = 8'hfa;
     14'b01010100111110: fc_kernel = 8'h02;
     14'b01010100111111: fc_kernel = 8'h04;
     14'b01010101000000: fc_kernel = 8'h0a;
     14'b01010101000001: fc_kernel = 8'h0b;
     14'b01010101000010: fc_kernel = 8'h08;
     14'b01010101000011: fc_kernel = 8'h03;
     14'b01010101000100: fc_kernel = 8'hf9;
     14'b01010101000101: fc_kernel = 8'hef;
     14'b01010101000110: fc_kernel = 8'heb;
     14'b01010101000111: fc_kernel = 8'hf6;
     14'b01010101001000: fc_kernel = 8'hf6;
     14'b01010101001001: fc_kernel = 8'hff;
     14'b01010101001010: fc_kernel = 8'hf5;
     14'b01010101001011: fc_kernel = 8'hfb;
     14'b01010101001100: fc_kernel = 8'hfc;
     14'b01010101001101: fc_kernel = 8'h06;
     14'b01010101001110: fc_kernel = 8'hff;
     14'b01010101001111: fc_kernel = 8'hed;
     14'b01010101010000: fc_kernel = 8'h07;
     14'b01010101010001: fc_kernel = 8'h01;
     14'b01010101010010: fc_kernel = 8'hfe;
     14'b01010101010011: fc_kernel = 8'hf9;
     14'b01010101010100: fc_kernel = 8'hf1;
     14'b01010101010101: fc_kernel = 8'hed;
     14'b01010101010110: fc_kernel = 8'hf3;
     14'b01010101010111: fc_kernel = 8'hfe;
     14'b01010101011000: fc_kernel = 8'h00;
     14'b01010101011001: fc_kernel = 8'h03;
     14'b01010101011010: fc_kernel = 8'h00;
     14'b01010101011011: fc_kernel = 8'hf8;
     14'b01010101011100: fc_kernel = 8'hef;
     14'b01010101011101: fc_kernel = 8'hee;
     14'b01010101011110: fc_kernel = 8'hf1;
     14'b01010101011111: fc_kernel = 8'hf8;
     14'b01010101100000: fc_kernel = 8'hfc;
     14'b01010101100001: fc_kernel = 8'h03;
     14'b01010101100010: fc_kernel = 8'hfe;
     14'b01010101100011: fc_kernel = 8'h00;
     14'b01010101100100: fc_kernel = 8'hfe;
     14'b01010101100101: fc_kernel = 8'h03;
     14'b01010101100110: fc_kernel = 8'h0a;
     14'b01010101100111: fc_kernel = 8'hf6;
     14'b01010101101000: fc_kernel = 8'h08;
     14'b01010101101001: fc_kernel = 8'hfd;
     14'b01010101101010: fc_kernel = 8'h03;
     14'b01010101101011: fc_kernel = 8'h0d;
     14'b01010101101100: fc_kernel = 8'h06;
     14'b01010101101101: fc_kernel = 8'hf9;
     14'b01010101101110: fc_kernel = 8'hf0;
     14'b01010101101111: fc_kernel = 8'hf0;
     14'b01010101110000: fc_kernel = 8'hf1;
     14'b01010101110001: fc_kernel = 8'hf8;
     14'b01010101110010: fc_kernel = 8'hf1;
     14'b01010101110011: fc_kernel = 8'he9;
     14'b01010101110100: fc_kernel = 8'hee;
     14'b01010101110101: fc_kernel = 8'hf4;
     14'b01010101110110: fc_kernel = 8'hfb;
     14'b01010101110111: fc_kernel = 8'hfe;
     14'b01010101111000: fc_kernel = 8'hfe;
     14'b01010101111001: fc_kernel = 8'h00;
     14'b01010101111010: fc_kernel = 8'hff;
     14'b01010101111011: fc_kernel = 8'hfd;
     14'b01010101111100: fc_kernel = 8'h01;
     14'b01010101111101: fc_kernel = 8'h02;
     14'b01010101111110: fc_kernel = 8'h0a;
     14'b01010101111111: fc_kernel = 8'hf3;
     14'b01010110000000: fc_kernel = 8'hf5;
     14'b01010110000001: fc_kernel = 8'h05;
     14'b01010110000010: fc_kernel = 8'h04;
     14'b01010110000011: fc_kernel = 8'h09;
     14'b01010110000100: fc_kernel = 8'h0b;
     14'b01010110000101: fc_kernel = 8'h06;
     14'b01010110000110: fc_kernel = 8'hf6;
     14'b01010110000111: fc_kernel = 8'hf3;
     14'b01010110001000: fc_kernel = 8'hf4;
     14'b01010110001001: fc_kernel = 8'hfa;
     14'b01010110001010: fc_kernel = 8'hf5;
     14'b01010110001011: fc_kernel = 8'hf3;
     14'b01010110001100: fc_kernel = 8'hfc;
     14'b01010110001101: fc_kernel = 8'hfb;
     14'b01010110001110: fc_kernel = 8'hff;
     14'b01010110001111: fc_kernel = 8'h01;
     14'b01010110010000: fc_kernel = 8'h01;
     14'b01010110010001: fc_kernel = 8'hfe;
     14'b01010110010010: fc_kernel = 8'h05;
     14'b01010110010011: fc_kernel = 8'h01;
     14'b01010110010100: fc_kernel = 8'hff;
     14'b01010110010101: fc_kernel = 8'h05;
     14'b01010110010110: fc_kernel = 8'h05;
     14'b01010110010111: fc_kernel = 8'hfd;
     14'b01010110011000: fc_kernel = 8'h12;
     14'b01010110011001: fc_kernel = 8'h09;
     14'b01010110011010: fc_kernel = 8'h04;
     14'b01010110011011: fc_kernel = 8'h03;
     14'b01010110011100: fc_kernel = 8'h02;
     14'b01010110011101: fc_kernel = 8'h02;
     14'b01010110011110: fc_kernel = 8'h01;
     14'b01010110011111: fc_kernel = 8'hfe;
     14'b01010110100000: fc_kernel = 8'hfa;
     14'b01010110100001: fc_kernel = 8'hf9;
     14'b01010110100010: fc_kernel = 8'hf9;
     14'b01010110100011: fc_kernel = 8'hf7;
     14'b01010110100100: fc_kernel = 8'hff;
     14'b01010110100101: fc_kernel = 8'hf8;
     14'b01010110100110: fc_kernel = 8'hfe;
     14'b01010110100111: fc_kernel = 8'h01;
     14'b01010110101000: fc_kernel = 8'h00;
     14'b01010110101001: fc_kernel = 8'h02;
     14'b01010110101010: fc_kernel = 8'h02;
     14'b01010110101011: fc_kernel = 8'h03;
     14'b01010110101100: fc_kernel = 8'h02;
     14'b01010110101101: fc_kernel = 8'h09;
     14'b01010110101110: fc_kernel = 8'h06;
     14'b01010110101111: fc_kernel = 8'hfd;
     14'b01010110110000: fc_kernel = 8'h18;
     14'b01010110110001: fc_kernel = 8'h07;
     14'b01010110110010: fc_kernel = 8'h02;
     14'b01010110110011: fc_kernel = 8'h08;
     14'b01010110110100: fc_kernel = 8'h02;
     14'b01010110110101: fc_kernel = 8'h00;
     14'b01010110110110: fc_kernel = 8'h00;
     14'b01010110110111: fc_kernel = 8'h00;
     14'b01010110111000: fc_kernel = 8'h00;
     14'b01010110111001: fc_kernel = 8'h00;
     14'b01010110111010: fc_kernel = 8'h00;
     14'b01010110111011: fc_kernel = 8'hf7;
     14'b01010110111100: fc_kernel = 8'hfb;
     14'b01010110111101: fc_kernel = 8'h00;
     14'b01010110111110: fc_kernel = 8'h00;
     14'b01010110111111: fc_kernel = 8'h02;
     14'b01010111000000: fc_kernel = 8'h00;
     14'b01010111000001: fc_kernel = 8'hff;
     14'b01010111000010: fc_kernel = 8'hff;
     14'b01010111000011: fc_kernel = 8'h00;
     14'b01010111000100: fc_kernel = 8'h04;
     14'b01010111000101: fc_kernel = 8'h0d;
     14'b01010111000110: fc_kernel = 8'h01;
     14'b01010111000111: fc_kernel = 8'hf6;
     14'b01010111001000: fc_kernel = 8'h02;
     14'b01010111001001: fc_kernel = 8'h05;
     14'b01010111001010: fc_kernel = 8'h02;
     14'b01010111001011: fc_kernel = 8'hfd;
     14'b01010111001100: fc_kernel = 8'hfd;
     14'b01010111001101: fc_kernel = 8'hfe;
     14'b01010111001110: fc_kernel = 8'h00;
     14'b01010111001111: fc_kernel = 8'h01;
     14'b01010111010000: fc_kernel = 8'hfb;
     14'b01010111010001: fc_kernel = 8'h00;
     14'b01010111010010: fc_kernel = 8'h04;
     14'b01010111010011: fc_kernel = 8'hff;
     14'b01010111010100: fc_kernel = 8'h00;
     14'b01010111010101: fc_kernel = 8'hfd;
     14'b01010111010110: fc_kernel = 8'h04;
     14'b01010111010111: fc_kernel = 8'h04;
     14'b01010111011000: fc_kernel = 8'h04;
     14'b01010111011001: fc_kernel = 8'h07;
     14'b01010111011010: fc_kernel = 8'h02;
     14'b01010111011011: fc_kernel = 8'h08;
     14'b01010111011100: fc_kernel = 8'h08;
     14'b01010111011101: fc_kernel = 8'h08;
     14'b01010111011110: fc_kernel = 8'h05;
     14'b01010111011111: fc_kernel = 8'h03;
     14'b01010111100000: fc_kernel = 8'hf8;
     14'b01010111100001: fc_kernel = 8'h02;
     14'b01010111100010: fc_kernel = 8'h00;
     14'b01010111100011: fc_kernel = 8'hff;
     14'b01010111100100: fc_kernel = 8'hf7;
     14'b01010111100101: fc_kernel = 8'hfb;
     14'b01010111100110: fc_kernel = 8'h00;
     14'b01010111100111: fc_kernel = 8'hfc;
     14'b01010111101000: fc_kernel = 8'h00;
     14'b01010111101001: fc_kernel = 8'hfe;
     14'b01010111101010: fc_kernel = 8'h01;
     14'b01010111101011: fc_kernel = 8'h05;
     14'b01010111101100: fc_kernel = 8'hff;
     14'b01010111101101: fc_kernel = 8'h04;
     14'b01010111101110: fc_kernel = 8'h01;
     14'b01010111101111: fc_kernel = 8'h06;
     14'b01010111110000: fc_kernel = 8'h00;
     14'b01010111110001: fc_kernel = 8'h00;
     14'b01010111110010: fc_kernel = 8'h07;
     14'b01010111110011: fc_kernel = 8'h07;
     14'b01010111110100: fc_kernel = 8'h01;
     14'b01010111110101: fc_kernel = 8'h02;
     14'b01010111110110: fc_kernel = 8'h0a;
     14'b01010111110111: fc_kernel = 8'h09;
     14'b01010111111000: fc_kernel = 8'h04;
     14'b01010111111001: fc_kernel = 8'h03;
     14'b01010111111010: fc_kernel = 8'h0b;
     14'b01010111111011: fc_kernel = 8'h01;
     14'b01010111111100: fc_kernel = 8'hfb;
     14'b01010111111101: fc_kernel = 8'hfb;
     14'b01010111111110: fc_kernel = 8'hff;
     14'b01010111111111: fc_kernel = 8'h02;
     14'b01011000000000: fc_kernel = 8'h02;
     14'b01011000000001: fc_kernel = 8'h02;
     14'b01011000000010: fc_kernel = 8'h04;
     14'b01011000000011: fc_kernel = 8'h01;
     14'b01011000000100: fc_kernel = 8'h01;
     14'b01011000000101: fc_kernel = 8'h05;
     14'b01011000000110: fc_kernel = 8'h02;
     14'b01011000000111: fc_kernel = 8'h00;
     14'b01011000001000: fc_kernel = 8'hfe;
     14'b01011000001001: fc_kernel = 8'h02;
     14'b01011000001010: fc_kernel = 8'h00;
     14'b01011000001011: fc_kernel = 8'hff;
     14'b01011000001100: fc_kernel = 8'hfd;
     14'b01011000001101: fc_kernel = 8'h00;
     14'b01011000001110: fc_kernel = 8'h06;
     14'b01011000001111: fc_kernel = 8'h01;
     14'b01011000010000: fc_kernel = 8'h17;
     14'b01011000010001: fc_kernel = 8'h0d;
     14'b01011000010010: fc_kernel = 8'h03;
     14'b01011000010011: fc_kernel = 8'h06;
     14'b01011000010100: fc_kernel = 8'hff;
     14'b01011000010101: fc_kernel = 8'hf9;
     14'b01011000010110: fc_kernel = 8'h00;
     14'b01011000010111: fc_kernel = 8'h02;
     14'b01011000011000: fc_kernel = 8'h02;
     14'b01011000011001: fc_kernel = 8'h03;
     14'b01011000011010: fc_kernel = 8'h03;
     14'b01011000011011: fc_kernel = 8'h0a;
     14'b01011000011100: fc_kernel = 8'h03;
     14'b01011000011101: fc_kernel = 8'h08;
     14'b01011000011110: fc_kernel = 8'h05;
     14'b01011000011111: fc_kernel = 8'h07;
     14'b01011000100000: fc_kernel = 8'h01;
     14'b01011000100001: fc_kernel = 8'h00;
     14'b01011000100010: fc_kernel = 8'hff;
     14'b01011000100011: fc_kernel = 8'h06;
     14'b01011000100100: fc_kernel = 8'h0a;
     14'b01011000100101: fc_kernel = 8'h11;
     14'b01011000100110: fc_kernel = 8'h10;
     14'b01011000100111: fc_kernel = 8'h07;
     14'b01011000101000: fc_kernel = 8'h17;
     14'b01011000101001: fc_kernel = 8'h1d;
     14'b01011000101010: fc_kernel = 8'h10;
     14'b01011000101011: fc_kernel = 8'hfe;
     14'b01011000101100: fc_kernel = 8'hfb;
     14'b01011000101101: fc_kernel = 8'hf8;
     14'b01011000101110: fc_kernel = 8'h00;
     14'b01011000101111: fc_kernel = 8'h02;
     14'b01011000110000: fc_kernel = 8'h0b;
     14'b01011000110001: fc_kernel = 8'h02;
     14'b01011000110010: fc_kernel = 8'h0c;
     14'b01011000110011: fc_kernel = 8'h0c;
     14'b01011000110100: fc_kernel = 8'h0d;
     14'b01011000110101: fc_kernel = 8'h0b;
     14'b01011000110110: fc_kernel = 8'h10;
     14'b01011000110111: fc_kernel = 8'h11;
     14'b01011000111000: fc_kernel = 8'h0e;
     14'b01011000111001: fc_kernel = 8'h0d;
     14'b01011000111010: fc_kernel = 8'h0e;
     14'b01011000111011: fc_kernel = 8'h12;
     14'b01011000111100: fc_kernel = 8'h1f;
     14'b01011000111101: fc_kernel = 8'h24;
     14'b01011000111110: fc_kernel = 8'h18;
     14'b01011000111111: fc_kernel = 8'h0d;
     14'b01100000000000: fc_kernel = 8'h10;
     14'b01100000000001: fc_kernel = 8'h02;
     14'b01100000000010: fc_kernel = 8'hfe;
     14'b01100000000011: fc_kernel = 8'h02;
     14'b01100000000100: fc_kernel = 8'h31;
     14'b01100000000101: fc_kernel = 8'h1f;
     14'b01100000000110: fc_kernel = 8'h25;
     14'b01100000000111: fc_kernel = 8'h21;
     14'b01100000001000: fc_kernel = 8'h1f;
     14'b01100000001001: fc_kernel = 8'h1f;
     14'b01100000001010: fc_kernel = 8'h15;
     14'b01100000001011: fc_kernel = 8'h12;
     14'b01100000001100: fc_kernel = 8'h0f;
     14'b01100000001101: fc_kernel = 8'h09;
     14'b01100000001110: fc_kernel = 8'h07;
     14'b01100000001111: fc_kernel = 8'h0a;
     14'b01100000010000: fc_kernel = 8'h11;
     14'b01100000010001: fc_kernel = 8'h1d;
     14'b01100000010010: fc_kernel = 8'h1e;
     14'b01100000010011: fc_kernel = 8'h24;
     14'b01100000010100: fc_kernel = 8'h26;
     14'b01100000010101: fc_kernel = 8'h21;
     14'b01100000010110: fc_kernel = 8'h0a;
     14'b01100000010111: fc_kernel = 8'hfc;
     14'b01100000011000: fc_kernel = 8'h15;
     14'b01100000011001: fc_kernel = 8'heb;
     14'b01100000011010: fc_kernel = 8'h15;
     14'b01100000011011: fc_kernel = 8'h18;
     14'b01100000011100: fc_kernel = 8'h13;
     14'b01100000011101: fc_kernel = 8'h13;
     14'b01100000011110: fc_kernel = 8'h09;
     14'b01100000011111: fc_kernel = 8'h0c;
     14'b01100000100000: fc_kernel = 8'h09;
     14'b01100000100001: fc_kernel = 8'h06;
     14'b01100000100010: fc_kernel = 8'h04;
     14'b01100000100011: fc_kernel = 8'hff;
     14'b01100000100100: fc_kernel = 8'h00;
     14'b01100000100101: fc_kernel = 8'h01;
     14'b01100000100110: fc_kernel = 8'hfd;
     14'b01100000100111: fc_kernel = 8'hfe;
     14'b01100000101000: fc_kernel = 8'h01;
     14'b01100000101001: fc_kernel = 8'h01;
     14'b01100000101010: fc_kernel = 8'hfd;
     14'b01100000101011: fc_kernel = 8'h05;
     14'b01100000101100: fc_kernel = 8'h10;
     14'b01100000101101: fc_kernel = 8'h13;
     14'b01100000101110: fc_kernel = 8'h0b;
     14'b01100000101111: fc_kernel = 8'hff;
     14'b01100000110000: fc_kernel = 8'hfc;
     14'b01100000110001: fc_kernel = 8'hef;
     14'b01100000110010: fc_kernel = 8'h00;
     14'b01100000110011: fc_kernel = 8'h0c;
     14'b01100000110100: fc_kernel = 8'h01;
     14'b01100000110101: fc_kernel = 8'hfb;
     14'b01100000110110: fc_kernel = 8'hfd;
     14'b01100000110111: fc_kernel = 8'h03;
     14'b01100000111000: fc_kernel = 8'hfb;
     14'b01100000111001: fc_kernel = 8'hfa;
     14'b01100000111010: fc_kernel = 8'hf8;
     14'b01100000111011: fc_kernel = 8'hfc;
     14'b01100000111100: fc_kernel = 8'hfb;
     14'b01100000111101: fc_kernel = 8'hfc;
     14'b01100000111110: fc_kernel = 8'hf8;
     14'b01100000111111: fc_kernel = 8'hfb;
     14'b01100001000000: fc_kernel = 8'h03;
     14'b01100001000001: fc_kernel = 8'h00;
     14'b01100001000010: fc_kernel = 8'h06;
     14'b01100001000011: fc_kernel = 8'h03;
     14'b01100001000100: fc_kernel = 8'h0b;
     14'b01100001000101: fc_kernel = 8'h0b;
     14'b01100001000110: fc_kernel = 8'hfd;
     14'b01100001000111: fc_kernel = 8'hf5;
     14'b01100001001000: fc_kernel = 8'heb;
     14'b01100001001001: fc_kernel = 8'hf5;
     14'b01100001001010: fc_kernel = 8'hf7;
     14'b01100001001011: fc_kernel = 8'hf8;
     14'b01100001001100: fc_kernel = 8'hf6;
     14'b01100001001101: fc_kernel = 8'hf8;
     14'b01100001001110: fc_kernel = 8'hfa;
     14'b01100001001111: fc_kernel = 8'h01;
     14'b01100001010000: fc_kernel = 8'hfa;
     14'b01100001010001: fc_kernel = 8'hef;
     14'b01100001010010: fc_kernel = 8'hf2;
     14'b01100001010011: fc_kernel = 8'hf3;
     14'b01100001010100: fc_kernel = 8'hf4;
     14'b01100001010101: fc_kernel = 8'hf6;
     14'b01100001010110: fc_kernel = 8'hf8;
     14'b01100001010111: fc_kernel = 8'h01;
     14'b01100001011000: fc_kernel = 8'h02;
     14'b01100001011001: fc_kernel = 8'h04;
     14'b01100001011010: fc_kernel = 8'h06;
     14'b01100001011011: fc_kernel = 8'h04;
     14'b01100001011100: fc_kernel = 8'h08;
     14'b01100001011101: fc_kernel = 8'h0d;
     14'b01100001011110: fc_kernel = 8'h04;
     14'b01100001011111: fc_kernel = 8'hfa;
     14'b01100001100000: fc_kernel = 8'hd4;
     14'b01100001100001: fc_kernel = 8'hf1;
     14'b01100001100010: fc_kernel = 8'hf7;
     14'b01100001100011: fc_kernel = 8'hf3;
     14'b01100001100100: fc_kernel = 8'hed;
     14'b01100001100101: fc_kernel = 8'hf4;
     14'b01100001100110: fc_kernel = 8'hf9;
     14'b01100001100111: fc_kernel = 8'hf5;
     14'b01100001101000: fc_kernel = 8'hed;
     14'b01100001101001: fc_kernel = 8'hef;
     14'b01100001101010: fc_kernel = 8'hea;
     14'b01100001101011: fc_kernel = 8'hf4;
     14'b01100001101100: fc_kernel = 8'hf5;
     14'b01100001101101: fc_kernel = 8'hfb;
     14'b01100001101110: fc_kernel = 8'hf6;
     14'b01100001101111: fc_kernel = 8'hf8;
     14'b01100001110000: fc_kernel = 8'hfc;
     14'b01100001110001: fc_kernel = 8'h01;
     14'b01100001110010: fc_kernel = 8'h03;
     14'b01100001110011: fc_kernel = 8'h00;
     14'b01100001110100: fc_kernel = 8'h06;
     14'b01100001110101: fc_kernel = 8'h05;
     14'b01100001110110: fc_kernel = 8'h08;
     14'b01100001110111: fc_kernel = 8'h05;
     14'b01100001111000: fc_kernel = 8'hd9;
     14'b01100001111001: fc_kernel = 8'hec;
     14'b01100001111010: fc_kernel = 8'hf5;
     14'b01100001111011: fc_kernel = 8'hf9;
     14'b01100001111100: fc_kernel = 8'hef;
     14'b01100001111101: fc_kernel = 8'hf9;
     14'b01100001111110: fc_kernel = 8'hfd;
     14'b01100001111111: fc_kernel = 8'hf8;
     14'b01100010000000: fc_kernel = 8'hf8;
     14'b01100010000001: fc_kernel = 8'hfc;
     14'b01100010000010: fc_kernel = 8'hf7;
     14'b01100010000011: fc_kernel = 8'hf5;
     14'b01100010000100: fc_kernel = 8'hf6;
     14'b01100010000101: fc_kernel = 8'hf5;
     14'b01100010000110: fc_kernel = 8'hf8;
     14'b01100010000111: fc_kernel = 8'hf5;
     14'b01100010001000: fc_kernel = 8'hf4;
     14'b01100010001001: fc_kernel = 8'hf2;
     14'b01100010001010: fc_kernel = 8'hf8;
     14'b01100010001011: fc_kernel = 8'hfa;
     14'b01100010001100: fc_kernel = 8'hfc;
     14'b01100010001101: fc_kernel = 8'hfe;
     14'b01100010001110: fc_kernel = 8'h06;
     14'b01100010001111: fc_kernel = 8'h00;
     14'b01100010010000: fc_kernel = 8'hd1;
     14'b01100010010001: fc_kernel = 8'hfc;
     14'b01100010010010: fc_kernel = 8'hfc;
     14'b01100010010011: fc_kernel = 8'hf8;
     14'b01100010010100: fc_kernel = 8'hf1;
     14'b01100010010101: fc_kernel = 8'hf9;
     14'b01100010010110: fc_kernel = 8'hf6;
     14'b01100010010111: fc_kernel = 8'hee;
     14'b01100010011000: fc_kernel = 8'hf0;
     14'b01100010011001: fc_kernel = 8'hfc;
     14'b01100010011010: fc_kernel = 8'hf4;
     14'b01100010011011: fc_kernel = 8'hf1;
     14'b01100010011100: fc_kernel = 8'hf5;
     14'b01100010011101: fc_kernel = 8'hf2;
     14'b01100010011110: fc_kernel = 8'hf3;
     14'b01100010011111: fc_kernel = 8'hed;
     14'b01100010100000: fc_kernel = 8'hf0;
     14'b01100010100001: fc_kernel = 8'hed;
     14'b01100010100010: fc_kernel = 8'hf1;
     14'b01100010100011: fc_kernel = 8'hf4;
     14'b01100010100100: fc_kernel = 8'hf0;
     14'b01100010100101: fc_kernel = 8'hec;
     14'b01100010100110: fc_kernel = 8'hed;
     14'b01100010100111: fc_kernel = 8'hec;
     14'b01100010101000: fc_kernel = 8'hcf;
     14'b01100010101001: fc_kernel = 8'hfc;
     14'b01100010101010: fc_kernel = 8'hfa;
     14'b01100010101011: fc_kernel = 8'hef;
     14'b01100010101100: fc_kernel = 8'hee;
     14'b01100010101101: fc_kernel = 8'hf8;
     14'b01100010101110: fc_kernel = 8'hf7;
     14'b01100010101111: fc_kernel = 8'hf0;
     14'b01100010110000: fc_kernel = 8'hf3;
     14'b01100010110001: fc_kernel = 8'hf5;
     14'b01100010110010: fc_kernel = 8'hf5;
     14'b01100010110011: fc_kernel = 8'hee;
     14'b01100010110100: fc_kernel = 8'hf3;
     14'b01100010110101: fc_kernel = 8'heb;
     14'b01100010110110: fc_kernel = 8'he8;
     14'b01100010110111: fc_kernel = 8'he7;
     14'b01100010111000: fc_kernel = 8'he5;
     14'b01100010111001: fc_kernel = 8'he7;
     14'b01100010111010: fc_kernel = 8'hf4;
     14'b01100010111011: fc_kernel = 8'hf3;
     14'b01100010111100: fc_kernel = 8'heb;
     14'b01100010111101: fc_kernel = 8'he7;
     14'b01100010111110: fc_kernel = 8'hdb;
     14'b01100010111111: fc_kernel = 8'hc6;
     14'b01100011000000: fc_kernel = 8'hcf;
     14'b01100011000001: fc_kernel = 8'hf4;
     14'b01100011000010: fc_kernel = 8'hf8;
     14'b01100011000011: fc_kernel = 8'hea;
     14'b01100011000100: fc_kernel = 8'hef;
     14'b01100011000101: fc_kernel = 8'hf6;
     14'b01100011000110: fc_kernel = 8'hf7;
     14'b01100011000111: fc_kernel = 8'hf3;
     14'b01100011001000: fc_kernel = 8'hf6;
     14'b01100011001001: fc_kernel = 8'hf0;
     14'b01100011001010: fc_kernel = 8'hf2;
     14'b01100011001011: fc_kernel = 8'hf3;
     14'b01100011001100: fc_kernel = 8'hf0;
     14'b01100011001101: fc_kernel = 8'hea;
     14'b01100011001110: fc_kernel = 8'he7;
     14'b01100011001111: fc_kernel = 8'he5;
     14'b01100011010000: fc_kernel = 8'he5;
     14'b01100011010001: fc_kernel = 8'hf1;
     14'b01100011010010: fc_kernel = 8'hf5;
     14'b01100011010011: fc_kernel = 8'hf8;
     14'b01100011010100: fc_kernel = 8'hec;
     14'b01100011010101: fc_kernel = 8'hef;
     14'b01100011010110: fc_kernel = 8'hee;
     14'b01100011010111: fc_kernel = 8'hca;
     14'b01100011011000: fc_kernel = 8'hcb;
     14'b01100011011001: fc_kernel = 8'hf2;
     14'b01100011011010: fc_kernel = 8'hf1;
     14'b01100011011011: fc_kernel = 8'hec;
     14'b01100011011100: fc_kernel = 8'hf3;
     14'b01100011011101: fc_kernel = 8'hfe;
     14'b01100011011110: fc_kernel = 8'h00;
     14'b01100011011111: fc_kernel = 8'h00;
     14'b01100011100000: fc_kernel = 8'hfb;
     14'b01100011100001: fc_kernel = 8'hfd;
     14'b01100011100010: fc_kernel = 8'hfa;
     14'b01100011100011: fc_kernel = 8'hfb;
     14'b01100011100100: fc_kernel = 8'hf0;
     14'b01100011100101: fc_kernel = 8'he5;
     14'b01100011100110: fc_kernel = 8'heb;
     14'b01100011100111: fc_kernel = 8'hf0;
     14'b01100011101000: fc_kernel = 8'hf1;
     14'b01100011101001: fc_kernel = 8'hf7;
     14'b01100011101010: fc_kernel = 8'hfd;
     14'b01100011101011: fc_kernel = 8'hff;
     14'b01100011101100: fc_kernel = 8'hff;
     14'b01100011101101: fc_kernel = 8'h02;
     14'b01100011101110: fc_kernel = 8'hf9;
     14'b01100011101111: fc_kernel = 8'hd6;
     14'b01100011110000: fc_kernel = 8'hc7;
     14'b01100011110001: fc_kernel = 8'hf6;
     14'b01100011110010: fc_kernel = 8'hf7;
     14'b01100011110011: fc_kernel = 8'h00;
     14'b01100011110100: fc_kernel = 8'h00;
     14'b01100011110101: fc_kernel = 8'hff;
     14'b01100011110110: fc_kernel = 8'h02;
     14'b01100011110111: fc_kernel = 8'h03;
     14'b01100011111000: fc_kernel = 8'h00;
     14'b01100011111001: fc_kernel = 8'hfc;
     14'b01100011111010: fc_kernel = 8'h05;
     14'b01100011111011: fc_kernel = 8'h01;
     14'b01100011111100: fc_kernel = 8'hf4;
     14'b01100011111101: fc_kernel = 8'he8;
     14'b01100011111110: fc_kernel = 8'hf4;
     14'b01100011111111: fc_kernel = 8'hfa;
     14'b01100100000000: fc_kernel = 8'hf0;
     14'b01100100000001: fc_kernel = 8'hf7;
     14'b01100100000010: fc_kernel = 8'hf8;
     14'b01100100000011: fc_kernel = 8'h01;
     14'b01100100000100: fc_kernel = 8'h0b;
     14'b01100100000101: fc_kernel = 8'h1b;
     14'b01100100000110: fc_kernel = 8'h0f;
     14'b01100100000111: fc_kernel = 8'he7;
     14'b01100100001000: fc_kernel = 8'hcc;
     14'b01100100001001: fc_kernel = 8'hed;
     14'b01100100001010: fc_kernel = 8'h01;
     14'b01100100001011: fc_kernel = 8'h01;
     14'b01100100001100: fc_kernel = 8'h03;
     14'b01100100001101: fc_kernel = 8'h05;
     14'b01100100001110: fc_kernel = 8'hff;
     14'b01100100001111: fc_kernel = 8'hff;
     14'b01100100010000: fc_kernel = 8'hfd;
     14'b01100100010001: fc_kernel = 8'h00;
     14'b01100100010010: fc_kernel = 8'h07;
     14'b01100100010011: fc_kernel = 8'hfa;
     14'b01100100010100: fc_kernel = 8'hf1;
     14'b01100100010101: fc_kernel = 8'hf2;
     14'b01100100010110: fc_kernel = 8'hf9;
     14'b01100100010111: fc_kernel = 8'hf9;
     14'b01100100011000: fc_kernel = 8'hf9;
     14'b01100100011001: fc_kernel = 8'hf9;
     14'b01100100011010: fc_kernel = 8'hfc;
     14'b01100100011011: fc_kernel = 8'h04;
     14'b01100100011100: fc_kernel = 8'h0c;
     14'b01100100011101: fc_kernel = 8'h20;
     14'b01100100011110: fc_kernel = 8'h14;
     14'b01100100011111: fc_kernel = 8'hef;
     14'b01100100100000: fc_kernel = 8'hdc;
     14'b01100100100001: fc_kernel = 8'hda;
     14'b01100100100010: fc_kernel = 8'hf2;
     14'b01100100100011: fc_kernel = 8'h00;
     14'b01100100100100: fc_kernel = 8'h03;
     14'b01100100100101: fc_kernel = 8'hfe;
     14'b01100100100110: fc_kernel = 8'hfd;
     14'b01100100100111: fc_kernel = 8'h05;
     14'b01100100101000: fc_kernel = 8'h07;
     14'b01100100101001: fc_kernel = 8'h07;
     14'b01100100101010: fc_kernel = 8'h00;
     14'b01100100101011: fc_kernel = 8'hfb;
     14'b01100100101100: fc_kernel = 8'hf6;
     14'b01100100101101: fc_kernel = 8'hfb;
     14'b01100100101110: fc_kernel = 8'h00;
     14'b01100100101111: fc_kernel = 8'hf4;
     14'b01100100110000: fc_kernel = 8'hf8;
     14'b01100100110001: fc_kernel = 8'h00;
     14'b01100100110010: fc_kernel = 8'hff;
     14'b01100100110011: fc_kernel = 8'h05;
     14'b01100100110100: fc_kernel = 8'h0a;
     14'b01100100110101: fc_kernel = 8'h1a;
     14'b01100100110110: fc_kernel = 8'h14;
     14'b01100100110111: fc_kernel = 8'hf5;
     14'b01100100111000: fc_kernel = 8'hd4;
     14'b01100100111001: fc_kernel = 8'hcc;
     14'b01100100111010: fc_kernel = 8'hf0;
     14'b01100100111011: fc_kernel = 8'h04;
     14'b01100100111100: fc_kernel = 8'h04;
     14'b01100100111101: fc_kernel = 8'h00;
     14'b01100100111110: fc_kernel = 8'h05;
     14'b01100100111111: fc_kernel = 8'h07;
     14'b01100101000000: fc_kernel = 8'h04;
     14'b01100101000001: fc_kernel = 8'h0e;
     14'b01100101000010: fc_kernel = 8'h04;
     14'b01100101000011: fc_kernel = 8'h00;
     14'b01100101000100: fc_kernel = 8'hfd;
     14'b01100101000101: fc_kernel = 8'h00;
     14'b01100101000110: fc_kernel = 8'h00;
     14'b01100101000111: fc_kernel = 8'hfb;
     14'b01100101001000: fc_kernel = 8'hf8;
     14'b01100101001001: fc_kernel = 8'hf9;
     14'b01100101001010: fc_kernel = 8'h03;
     14'b01100101001011: fc_kernel = 8'h03;
     14'b01100101001100: fc_kernel = 8'h03;
     14'b01100101001101: fc_kernel = 8'h04;
     14'b01100101001110: fc_kernel = 8'h03;
     14'b01100101001111: fc_kernel = 8'hf8;
     14'b01100101010000: fc_kernel = 8'hd7;
     14'b01100101010001: fc_kernel = 8'hba;
     14'b01100101010010: fc_kernel = 8'hee;
     14'b01100101010011: fc_kernel = 8'hfd;
     14'b01100101010100: fc_kernel = 8'h05;
     14'b01100101010101: fc_kernel = 8'h0c;
     14'b01100101010110: fc_kernel = 8'h08;
     14'b01100101010111: fc_kernel = 8'h08;
     14'b01100101011000: fc_kernel = 8'h14;
     14'b01100101011001: fc_kernel = 8'h11;
     14'b01100101011010: fc_kernel = 8'h07;
     14'b01100101011011: fc_kernel = 8'hfb;
     14'b01100101011100: fc_kernel = 8'h02;
     14'b01100101011101: fc_kernel = 8'hff;
     14'b01100101011110: fc_kernel = 8'hfb;
     14'b01100101011111: fc_kernel = 8'hf4;
     14'b01100101100000: fc_kernel = 8'hfe;
     14'b01100101100001: fc_kernel = 8'h04;
     14'b01100101100010: fc_kernel = 8'h02;
     14'b01100101100011: fc_kernel = 8'h05;
     14'b01100101100100: fc_kernel = 8'h03;
     14'b01100101100101: fc_kernel = 8'h00;
     14'b01100101100110: fc_kernel = 8'h00;
     14'b01100101100111: fc_kernel = 8'hfc;
     14'b01100101101000: fc_kernel = 8'hde;
     14'b01100101101001: fc_kernel = 8'hce;
     14'b01100101101010: fc_kernel = 8'hed;
     14'b01100101101011: fc_kernel = 8'hfa;
     14'b01100101101100: fc_kernel = 8'hff;
     14'b01100101101101: fc_kernel = 8'h09;
     14'b01100101101110: fc_kernel = 8'h09;
     14'b01100101101111: fc_kernel = 8'h0b;
     14'b01100101110000: fc_kernel = 8'h11;
     14'b01100101110001: fc_kernel = 8'h18;
     14'b01100101110010: fc_kernel = 8'h07;
     14'b01100101110011: fc_kernel = 8'hfe;
     14'b01100101110100: fc_kernel = 8'h03;
     14'b01100101110101: fc_kernel = 8'hff;
     14'b01100101110110: fc_kernel = 8'hf9;
     14'b01100101110111: fc_kernel = 8'hfc;
     14'b01100101111000: fc_kernel = 8'h02;
     14'b01100101111001: fc_kernel = 8'h06;
     14'b01100101111010: fc_kernel = 8'h03;
     14'b01100101111011: fc_kernel = 8'h06;
     14'b01100101111100: fc_kernel = 8'h06;
     14'b01100101111101: fc_kernel = 8'h02;
     14'b01100101111110: fc_kernel = 8'h09;
     14'b01100101111111: fc_kernel = 8'h00;
     14'b01100110000000: fc_kernel = 8'he5;
     14'b01100110000001: fc_kernel = 8'hdd;
     14'b01100110000010: fc_kernel = 8'hea;
     14'b01100110000011: fc_kernel = 8'hf8;
     14'b01100110000100: fc_kernel = 8'hfe;
     14'b01100110000101: fc_kernel = 8'h02;
     14'b01100110000110: fc_kernel = 8'h05;
     14'b01100110000111: fc_kernel = 8'h0d;
     14'b01100110001000: fc_kernel = 8'h15;
     14'b01100110001001: fc_kernel = 8'h17;
     14'b01100110001010: fc_kernel = 8'h10;
     14'b01100110001011: fc_kernel = 8'h07;
     14'b01100110001100: fc_kernel = 8'h04;
     14'b01100110001101: fc_kernel = 8'h00;
     14'b01100110001110: fc_kernel = 8'h03;
     14'b01100110001111: fc_kernel = 8'h05;
     14'b01100110010000: fc_kernel = 8'h07;
     14'b01100110010001: fc_kernel = 8'h07;
     14'b01100110010010: fc_kernel = 8'h02;
     14'b01100110010011: fc_kernel = 8'h04;
     14'b01100110010100: fc_kernel = 8'h01;
     14'b01100110010101: fc_kernel = 8'h00;
     14'b01100110010110: fc_kernel = 8'h07;
     14'b01100110010111: fc_kernel = 8'h03;
     14'b01100110011000: fc_kernel = 8'he2;
     14'b01100110011001: fc_kernel = 8'he9;
     14'b01100110011010: fc_kernel = 8'hee;
     14'b01100110011011: fc_kernel = 8'hf7;
     14'b01100110011100: fc_kernel = 8'hff;
     14'b01100110011101: fc_kernel = 8'hfe;
     14'b01100110011110: fc_kernel = 8'h06;
     14'b01100110011111: fc_kernel = 8'h07;
     14'b01100110100000: fc_kernel = 8'h0c;
     14'b01100110100001: fc_kernel = 8'h12;
     14'b01100110100010: fc_kernel = 8'h16;
     14'b01100110100011: fc_kernel = 8'h12;
     14'b01100110100100: fc_kernel = 8'h04;
     14'b01100110100101: fc_kernel = 8'h08;
     14'b01100110100110: fc_kernel = 8'h05;
     14'b01100110100111: fc_kernel = 8'h0a;
     14'b01100110101000: fc_kernel = 8'h08;
     14'b01100110101001: fc_kernel = 8'h00;
     14'b01100110101010: fc_kernel = 8'h05;
     14'b01100110101011: fc_kernel = 8'h05;
     14'b01100110101100: fc_kernel = 8'h02;
     14'b01100110101101: fc_kernel = 8'hfe;
     14'b01100110101110: fc_kernel = 8'h02;
     14'b01100110101111: fc_kernel = 8'hfa;
     14'b01100110110000: fc_kernel = 8'he6;
     14'b01100110110001: fc_kernel = 8'he5;
     14'b01100110110010: fc_kernel = 8'he6;
     14'b01100110110011: fc_kernel = 8'hf0;
     14'b01100110110100: fc_kernel = 8'hff;
     14'b01100110110101: fc_kernel = 8'h03;
     14'b01100110110110: fc_kernel = 8'h00;
     14'b01100110110111: fc_kernel = 8'h07;
     14'b01100110111000: fc_kernel = 8'h12;
     14'b01100110111001: fc_kernel = 8'h14;
     14'b01100110111010: fc_kernel = 8'h12;
     14'b01100110111011: fc_kernel = 8'h10;
     14'b01100110111100: fc_kernel = 8'h15;
     14'b01100110111101: fc_kernel = 8'h10;
     14'b01100110111110: fc_kernel = 8'h0f;
     14'b01100110111111: fc_kernel = 8'h07;
     14'b01100111000000: fc_kernel = 8'h0c;
     14'b01100111000001: fc_kernel = 8'h08;
     14'b01100111000010: fc_kernel = 8'h05;
     14'b01100111000011: fc_kernel = 8'h03;
     14'b01100111000100: fc_kernel = 8'h02;
     14'b01100111000101: fc_kernel = 8'h01;
     14'b01100111000110: fc_kernel = 8'h02;
     14'b01100111000111: fc_kernel = 8'hf9;
     14'b01100111001000: fc_kernel = 8'he5;
     14'b01100111001001: fc_kernel = 8'hdf;
     14'b01100111001010: fc_kernel = 8'he1;
     14'b01100111001011: fc_kernel = 8'he2;
     14'b01100111001100: fc_kernel = 8'hf0;
     14'b01100111001101: fc_kernel = 8'hfd;
     14'b01100111001110: fc_kernel = 8'h03;
     14'b01100111001111: fc_kernel = 8'h0a;
     14'b01100111010000: fc_kernel = 8'h10;
     14'b01100111010001: fc_kernel = 8'h16;
     14'b01100111010010: fc_kernel = 8'h12;
     14'b01100111010011: fc_kernel = 8'h13;
     14'b01100111010100: fc_kernel = 8'h10;
     14'b01100111010101: fc_kernel = 8'h08;
     14'b01100111010110: fc_kernel = 8'h08;
     14'b01100111010111: fc_kernel = 8'h0a;
     14'b01100111011000: fc_kernel = 8'h0a;
     14'b01100111011001: fc_kernel = 8'h04;
     14'b01100111011010: fc_kernel = 8'h02;
     14'b01100111011011: fc_kernel = 8'h02;
     14'b01100111011100: fc_kernel = 8'hfe;
     14'b01100111011101: fc_kernel = 8'hf6;
     14'b01100111011110: fc_kernel = 8'hf6;
     14'b01100111011111: fc_kernel = 8'hee;
     14'b01100111100000: fc_kernel = 8'he1;
     14'b01100111100001: fc_kernel = 8'hdd;
     14'b01100111100010: fc_kernel = 8'he1;
     14'b01100111100011: fc_kernel = 8'hd9;
     14'b01100111100100: fc_kernel = 8'he0;
     14'b01100111100101: fc_kernel = 8'hf4;
     14'b01100111100110: fc_kernel = 8'h02;
     14'b01100111100111: fc_kernel = 8'h0b;
     14'b01100111101000: fc_kernel = 8'h0b;
     14'b01100111101001: fc_kernel = 8'h0d;
     14'b01100111101010: fc_kernel = 8'h0c;
     14'b01100111101011: fc_kernel = 8'h0e;
     14'b01100111101100: fc_kernel = 8'h0f;
     14'b01100111101101: fc_kernel = 8'h0b;
     14'b01100111101110: fc_kernel = 8'h08;
     14'b01100111101111: fc_kernel = 8'h0a;
     14'b01100111110000: fc_kernel = 8'h06;
     14'b01100111110001: fc_kernel = 8'h08;
     14'b01100111110010: fc_kernel = 8'h01;
     14'b01100111110011: fc_kernel = 8'h02;
     14'b01100111110100: fc_kernel = 8'hfa;
     14'b01100111110101: fc_kernel = 8'hed;
     14'b01100111110110: fc_kernel = 8'he3;
     14'b01100111110111: fc_kernel = 8'he5;
     14'b01100111111000: fc_kernel = 8'he5;
     14'b01100111111001: fc_kernel = 8'he0;
     14'b01100111111010: fc_kernel = 8'hde;
     14'b01100111111011: fc_kernel = 8'hda;
     14'b01100111111100: fc_kernel = 8'hdf;
     14'b01100111111101: fc_kernel = 8'hec;
     14'b01100111111110: fc_kernel = 8'hf8;
     14'b01100111111111: fc_kernel = 8'h00;
     14'b01101000000000: fc_kernel = 8'hfd;
     14'b01101000000001: fc_kernel = 8'hff;
     14'b01101000000010: fc_kernel = 8'h04;
     14'b01101000000011: fc_kernel = 8'h01;
     14'b01101000000100: fc_kernel = 8'h03;
     14'b01101000000101: fc_kernel = 8'h01;
     14'b01101000000110: fc_kernel = 8'h07;
     14'b01101000000111: fc_kernel = 8'h00;
     14'b01101000001000: fc_kernel = 8'hfe;
     14'b01101000001001: fc_kernel = 8'h00;
     14'b01101000001010: fc_kernel = 8'h00;
     14'b01101000001011: fc_kernel = 8'h01;
     14'b01101000001100: fc_kernel = 8'hf5;
     14'b01101000001101: fc_kernel = 8'he5;
     14'b01101000001110: fc_kernel = 8'hdf;
     14'b01101000001111: fc_kernel = 8'he3;
     14'b01101000010000: fc_kernel = 8'he8;
     14'b01101000010001: fc_kernel = 8'he2;
     14'b01101000010010: fc_kernel = 8'hd2;
     14'b01101000010011: fc_kernel = 8'hca;
     14'b01101000010100: fc_kernel = 8'hdb;
     14'b01101000010101: fc_kernel = 8'hda;
     14'b01101000010110: fc_kernel = 8'hed;
     14'b01101000010111: fc_kernel = 8'he7;
     14'b01101000011000: fc_kernel = 8'he7;
     14'b01101000011001: fc_kernel = 8'he7;
     14'b01101000011010: fc_kernel = 8'hee;
     14'b01101000011011: fc_kernel = 8'hf5;
     14'b01101000011100: fc_kernel = 8'hf6;
     14'b01101000011101: fc_kernel = 8'hf5;
     14'b01101000011110: fc_kernel = 8'hf9;
     14'b01101000011111: fc_kernel = 8'hf5;
     14'b01101000100000: fc_kernel = 8'hfa;
     14'b01101000100001: fc_kernel = 8'hfd;
     14'b01101000100010: fc_kernel = 8'hfb;
     14'b01101000100011: fc_kernel = 8'hfa;
     14'b01101000100100: fc_kernel = 8'heb;
     14'b01101000100101: fc_kernel = 8'he4;
     14'b01101000100110: fc_kernel = 8'hdd;
     14'b01101000100111: fc_kernel = 8'he3;
     14'b01101000101000: fc_kernel = 8'hfa;
     14'b01101000101001: fc_kernel = 8'hf2;
     14'b01101000101010: fc_kernel = 8'he5;
     14'b01101000101011: fc_kernel = 8'hd5;
     14'b01101000101100: fc_kernel = 8'hd1;
     14'b01101000101101: fc_kernel = 8'hd6;
     14'b01101000101110: fc_kernel = 8'hdb;
     14'b01101000101111: fc_kernel = 8'hd3;
     14'b01101000110000: fc_kernel = 8'hc9;
     14'b01101000110001: fc_kernel = 8'hd9;
     14'b01101000110010: fc_kernel = 8'hea;
     14'b01101000110011: fc_kernel = 8'he5;
     14'b01101000110100: fc_kernel = 8'hd8;
     14'b01101000110101: fc_kernel = 8'hdd;
     14'b01101000110110: fc_kernel = 8'he8;
     14'b01101000110111: fc_kernel = 8'hef;
     14'b01101000111000: fc_kernel = 8'hed;
     14'b01101000111001: fc_kernel = 8'hea;
     14'b01101000111010: fc_kernel = 8'he3;
     14'b01101000111011: fc_kernel = 8'hea;
     14'b01101000111100: fc_kernel = 8'hdb;
     14'b01101000111101: fc_kernel = 8'hdb;
     14'b01101000111110: fc_kernel = 8'hdf;
     14'b01101000111111: fc_kernel = 8'he4;
     14'b01110000000000: fc_kernel = 8'hea;
     14'b01110000000001: fc_kernel = 8'he4;
     14'b01110000000010: fc_kernel = 8'hd0;
     14'b01110000000011: fc_kernel = 8'hd8;
     14'b01110000000100: fc_kernel = 8'hcf;
     14'b01110000000101: fc_kernel = 8'hcf;
     14'b01110000000110: fc_kernel = 8'hc5;
     14'b01110000000111: fc_kernel = 8'hec;
     14'b01110000001000: fc_kernel = 8'hcd;
     14'b01110000001001: fc_kernel = 8'hc8;
     14'b01110000001010: fc_kernel = 8'hcc;
     14'b01110000001011: fc_kernel = 8'hd5;
     14'b01110000001100: fc_kernel = 8'hd3;
     14'b01110000001101: fc_kernel = 8'hdd;
     14'b01110000001110: fc_kernel = 8'hdb;
     14'b01110000001111: fc_kernel = 8'he0;
     14'b01110000010000: fc_kernel = 8'he8;
     14'b01110000010001: fc_kernel = 8'hfc;
     14'b01110000010010: fc_kernel = 8'heb;
     14'b01110000010011: fc_kernel = 8'hf2;
     14'b01110000010100: fc_kernel = 8'hf4;
     14'b01110000010101: fc_kernel = 8'hf6;
     14'b01110000010110: fc_kernel = 8'hf0;
     14'b01110000010111: fc_kernel = 8'hf6;
     14'b01110000011000: fc_kernel = 8'he8;
     14'b01110000011001: fc_kernel = 8'h13;
     14'b01110000011010: fc_kernel = 8'hde;
     14'b01110000011011: fc_kernel = 8'hf4;
     14'b01110000011100: fc_kernel = 8'hfe;
     14'b01110000011101: fc_kernel = 8'hcd;
     14'b01110000011110: fc_kernel = 8'hc4;
     14'b01110000011111: fc_kernel = 8'hcf;
     14'b01110000100000: fc_kernel = 8'hd1;
     14'b01110000100001: fc_kernel = 8'hc8;
     14'b01110000100010: fc_kernel = 8'hd5;
     14'b01110000100011: fc_kernel = 8'hc4;
     14'b01110000100100: fc_kernel = 8'hcf;
     14'b01110000100101: fc_kernel = 8'hcc;
     14'b01110000100110: fc_kernel = 8'hc5;
     14'b01110000100111: fc_kernel = 8'hce;
     14'b01110000101000: fc_kernel = 8'hdc;
     14'b01110000101001: fc_kernel = 8'hed;
     14'b01110000101010: fc_kernel = 8'he2;
     14'b01110000101011: fc_kernel = 8'hdd;
     14'b01110000101100: fc_kernel = 8'hd4;
     14'b01110000101101: fc_kernel = 8'hdc;
     14'b01110000101110: fc_kernel = 8'he0;
     14'b01110000101111: fc_kernel = 8'hee;
     14'b01110000110000: fc_kernel = 8'hec;
     14'b01110000110001: fc_kernel = 8'h18;
     14'b01110000110010: fc_kernel = 8'hfc;
     14'b01110000110011: fc_kernel = 8'h04;
     14'b01110000110100: fc_kernel = 8'he6;
     14'b01110000110101: fc_kernel = 8'hfb;
     14'b01110000110110: fc_kernel = 8'h01;
     14'b01110000110111: fc_kernel = 8'heb;
     14'b01110000111000: fc_kernel = 8'hd4;
     14'b01110000111001: fc_kernel = 8'hd9;
     14'b01110000111010: fc_kernel = 8'hec;
     14'b01110000111011: fc_kernel = 8'he9;
     14'b01110000111100: fc_kernel = 8'he4;
     14'b01110000111101: fc_kernel = 8'hdc;
     14'b01110000111110: fc_kernel = 8'hda;
     14'b01110000111111: fc_kernel = 8'hd5;
     14'b01110001000000: fc_kernel = 8'hd7;
     14'b01110001000001: fc_kernel = 8'hd7;
     14'b01110001000010: fc_kernel = 8'he5;
     14'b01110001000011: fc_kernel = 8'he2;
     14'b01110001000100: fc_kernel = 8'hed;
     14'b01110001000101: fc_kernel = 8'hdf;
     14'b01110001000110: fc_kernel = 8'he6;
     14'b01110001000111: fc_kernel = 8'hec;
     14'b01110001001000: fc_kernel = 8'hf5;
     14'b01110001001001: fc_kernel = 8'h00;
     14'b01110001001010: fc_kernel = 8'h0f;
     14'b01110001001011: fc_kernel = 8'h18;
     14'b01110001001100: fc_kernel = 8'h16;
     14'b01110001001101: fc_kernel = 8'h1f;
     14'b01110001001110: fc_kernel = 8'h15;
     14'b01110001001111: fc_kernel = 8'h0f;
     14'b01110001010000: fc_kernel = 8'h0c;
     14'b01110001010001: fc_kernel = 8'h08;
     14'b01110001010010: fc_kernel = 8'h05;
     14'b01110001010011: fc_kernel = 8'h06;
     14'b01110001010100: fc_kernel = 8'h0a;
     14'b01110001010101: fc_kernel = 8'h00;
     14'b01110001010110: fc_kernel = 8'hfb;
     14'b01110001010111: fc_kernel = 8'hf5;
     14'b01110001011000: fc_kernel = 8'hf3;
     14'b01110001011001: fc_kernel = 8'he8;
     14'b01110001011010: fc_kernel = 8'hd7;
     14'b01110001011011: fc_kernel = 8'he0;
     14'b01110001011100: fc_kernel = 8'he2;
     14'b01110001011101: fc_kernel = 8'hda;
     14'b01110001011110: fc_kernel = 8'he0;
     14'b01110001011111: fc_kernel = 8'hee;
     14'b01110001100000: fc_kernel = 8'h1a;
     14'b01110001100001: fc_kernel = 8'h11;
     14'b01110001100010: fc_kernel = 8'h07;
     14'b01110001100011: fc_kernel = 8'h0c;
     14'b01110001100100: fc_kernel = 8'h0b;
     14'b01110001100101: fc_kernel = 8'h0c;
     14'b01110001100110: fc_kernel = 8'h0d;
     14'b01110001100111: fc_kernel = 8'h0e;
     14'b01110001101000: fc_kernel = 8'h0b;
     14'b01110001101001: fc_kernel = 8'h0b;
     14'b01110001101010: fc_kernel = 8'h0b;
     14'b01110001101011: fc_kernel = 8'h08;
     14'b01110001101100: fc_kernel = 8'hfd;
     14'b01110001101101: fc_kernel = 8'hfe;
     14'b01110001101110: fc_kernel = 8'h02;
     14'b01110001101111: fc_kernel = 8'h01;
     14'b01110001110000: fc_kernel = 8'hfc;
     14'b01110001110001: fc_kernel = 8'hf3;
     14'b01110001110010: fc_kernel = 8'hf9;
     14'b01110001110011: fc_kernel = 8'hfa;
     14'b01110001110100: fc_kernel = 8'hf8;
     14'b01110001110101: fc_kernel = 8'hef;
     14'b01110001110110: fc_kernel = 8'he6;
     14'b01110001110111: fc_kernel = 8'he3;
     14'b01110001111000: fc_kernel = 8'h2b;
     14'b01110001111001: fc_kernel = 8'h16;
     14'b01110001111010: fc_kernel = 8'h08;
     14'b01110001111011: fc_kernel = 8'h04;
     14'b01110001111100: fc_kernel = 8'h10;
     14'b01110001111101: fc_kernel = 8'h0f;
     14'b01110001111110: fc_kernel = 8'h0b;
     14'b01110001111111: fc_kernel = 8'h09;
     14'b01110010000000: fc_kernel = 8'h0b;
     14'b01110010000001: fc_kernel = 8'h0d;
     14'b01110010000010: fc_kernel = 8'h0c;
     14'b01110010000011: fc_kernel = 8'h07;
     14'b01110010000100: fc_kernel = 8'h00;
     14'b01110010000101: fc_kernel = 8'h07;
     14'b01110010000110: fc_kernel = 8'h06;
     14'b01110010000111: fc_kernel = 8'h09;
     14'b01110010001000: fc_kernel = 8'h08;
     14'b01110010001001: fc_kernel = 8'h05;
     14'b01110010001010: fc_kernel = 8'h05;
     14'b01110010001011: fc_kernel = 8'h00;
     14'b01110010001100: fc_kernel = 8'h00;
     14'b01110010001101: fc_kernel = 8'hf6;
     14'b01110010001110: fc_kernel = 8'hea;
     14'b01110010001111: fc_kernel = 8'he8;
     14'b01110010010000: fc_kernel = 8'h27;
     14'b01110010010001: fc_kernel = 8'h18;
     14'b01110010010010: fc_kernel = 8'h07;
     14'b01110010010011: fc_kernel = 8'h03;
     14'b01110010010100: fc_kernel = 8'h10;
     14'b01110010010101: fc_kernel = 8'h11;
     14'b01110010010110: fc_kernel = 8'h0f;
     14'b01110010010111: fc_kernel = 8'h08;
     14'b01110010011000: fc_kernel = 8'h10;
     14'b01110010011001: fc_kernel = 8'h11;
     14'b01110010011010: fc_kernel = 8'h13;
     14'b01110010011011: fc_kernel = 8'h0d;
     14'b01110010011100: fc_kernel = 8'h07;
     14'b01110010011101: fc_kernel = 8'h0c;
     14'b01110010011110: fc_kernel = 8'h10;
     14'b01110010011111: fc_kernel = 8'h0c;
     14'b01110010100000: fc_kernel = 8'h11;
     14'b01110010100001: fc_kernel = 8'h0d;
     14'b01110010100010: fc_kernel = 8'h02;
     14'b01110010100011: fc_kernel = 8'h01;
     14'b01110010100100: fc_kernel = 8'h00;
     14'b01110010100101: fc_kernel = 8'h07;
     14'b01110010100110: fc_kernel = 8'hf6;
     14'b01110010100111: fc_kernel = 8'he0;
     14'b01110010101000: fc_kernel = 8'h1d;
     14'b01110010101001: fc_kernel = 8'h10;
     14'b01110010101010: fc_kernel = 8'h09;
     14'b01110010101011: fc_kernel = 8'h06;
     14'b01110010101100: fc_kernel = 8'h0f;
     14'b01110010101101: fc_kernel = 8'h0e;
     14'b01110010101110: fc_kernel = 8'h0d;
     14'b01110010101111: fc_kernel = 8'h05;
     14'b01110010110000: fc_kernel = 8'h04;
     14'b01110010110001: fc_kernel = 8'h06;
     14'b01110010110010: fc_kernel = 8'h0e;
     14'b01110010110011: fc_kernel = 8'h09;
     14'b01110010110100: fc_kernel = 8'h0d;
     14'b01110010110101: fc_kernel = 8'h10;
     14'b01110010110110: fc_kernel = 8'h15;
     14'b01110010110111: fc_kernel = 8'h14;
     14'b01110010111000: fc_kernel = 8'h0f;
     14'b01110010111001: fc_kernel = 8'h0e;
     14'b01110010111010: fc_kernel = 8'h06;
     14'b01110010111011: fc_kernel = 8'h03;
     14'b01110010111100: fc_kernel = 8'h04;
     14'b01110010111101: fc_kernel = 8'hff;
     14'b01110010111110: fc_kernel = 8'hf4;
     14'b01110010111111: fc_kernel = 8'hee;
     14'b01110011000000: fc_kernel = 8'h1e;
     14'b01110011000001: fc_kernel = 8'h11;
     14'b01110011000010: fc_kernel = 8'h08;
     14'b01110011000011: fc_kernel = 8'h0d;
     14'b01110011000100: fc_kernel = 8'h0a;
     14'b01110011000101: fc_kernel = 8'h02;
     14'b01110011000110: fc_kernel = 8'hff;
     14'b01110011000111: fc_kernel = 8'h03;
     14'b01110011001000: fc_kernel = 8'h03;
     14'b01110011001001: fc_kernel = 8'h03;
     14'b01110011001010: fc_kernel = 8'h07;
     14'b01110011001011: fc_kernel = 8'h0c;
     14'b01110011001100: fc_kernel = 8'h0f;
     14'b01110011001101: fc_kernel = 8'h12;
     14'b01110011001110: fc_kernel = 8'h16;
     14'b01110011001111: fc_kernel = 8'h10;
     14'b01110011010000: fc_kernel = 8'h0d;
     14'b01110011010001: fc_kernel = 8'h0f;
     14'b01110011010010: fc_kernel = 8'h0a;
     14'b01110011010011: fc_kernel = 8'h0a;
     14'b01110011010100: fc_kernel = 8'h08;
     14'b01110011010101: fc_kernel = 8'hfc;
     14'b01110011010110: fc_kernel = 8'hf0;
     14'b01110011010111: fc_kernel = 8'hea;
     14'b01110011011000: fc_kernel = 8'h2a;
     14'b01110011011001: fc_kernel = 8'h13;
     14'b01110011011010: fc_kernel = 8'h07;
     14'b01110011011011: fc_kernel = 8'h03;
     14'b01110011011100: fc_kernel = 8'hff;
     14'b01110011011101: fc_kernel = 8'h00;
     14'b01110011011110: fc_kernel = 8'hff;
     14'b01110011011111: fc_kernel = 8'h03;
     14'b01110011100000: fc_kernel = 8'h04;
     14'b01110011100001: fc_kernel = 8'h02;
     14'b01110011100010: fc_kernel = 8'h02;
     14'b01110011100011: fc_kernel = 8'h08;
     14'b01110011100100: fc_kernel = 8'h12;
     14'b01110011100101: fc_kernel = 8'h17;
     14'b01110011100110: fc_kernel = 8'h19;
     14'b01110011100111: fc_kernel = 8'h17;
     14'b01110011101000: fc_kernel = 8'h14;
     14'b01110011101001: fc_kernel = 8'h11;
     14'b01110011101010: fc_kernel = 8'h0c;
     14'b01110011101011: fc_kernel = 8'h0e;
     14'b01110011101100: fc_kernel = 8'h07;
     14'b01110011101101: fc_kernel = 8'hfb;
     14'b01110011101110: fc_kernel = 8'he5;
     14'b01110011101111: fc_kernel = 8'he6;
     14'b01110011110000: fc_kernel = 8'h2d;
     14'b01110011110001: fc_kernel = 8'h21;
     14'b01110011110010: fc_kernel = 8'h0b;
     14'b01110011110011: fc_kernel = 8'h01;
     14'b01110011110100: fc_kernel = 8'h05;
     14'b01110011110101: fc_kernel = 8'h07;
     14'b01110011110110: fc_kernel = 8'h08;
     14'b01110011110111: fc_kernel = 8'h01;
     14'b01110011111000: fc_kernel = 8'h03;
     14'b01110011111001: fc_kernel = 8'hff;
     14'b01110011111010: fc_kernel = 8'hf4;
     14'b01110011111011: fc_kernel = 8'hea;
     14'b01110011111100: fc_kernel = 8'hfe;
     14'b01110011111101: fc_kernel = 8'h10;
     14'b01110011111110: fc_kernel = 8'h12;
     14'b01110011111111: fc_kernel = 8'h17;
     14'b01110100000000: fc_kernel = 8'h09;
     14'b01110100000001: fc_kernel = 8'h02;
     14'b01110100000010: fc_kernel = 8'h00;
     14'b01110100000011: fc_kernel = 8'h0a;
     14'b01110100000100: fc_kernel = 8'h02;
     14'b01110100000101: fc_kernel = 8'hef;
     14'b01110100000110: fc_kernel = 8'he8;
     14'b01110100000111: fc_kernel = 8'heb;
     14'b01110100001000: fc_kernel = 8'h2a;
     14'b01110100001001: fc_kernel = 8'h1f;
     14'b01110100001010: fc_kernel = 8'h13;
     14'b01110100001011: fc_kernel = 8'h07;
     14'b01110100001100: fc_kernel = 8'hff;
     14'b01110100001101: fc_kernel = 8'h09;
     14'b01110100001110: fc_kernel = 8'h04;
     14'b01110100001111: fc_kernel = 8'h02;
     14'b01110100010000: fc_kernel = 8'h03;
     14'b01110100010001: fc_kernel = 8'hf6;
     14'b01110100010010: fc_kernel = 8'hda;
     14'b01110100010011: fc_kernel = 8'hd3;
     14'b01110100010100: fc_kernel = 8'hf3;
     14'b01110100010101: fc_kernel = 8'h0b;
     14'b01110100010110: fc_kernel = 8'h10;
     14'b01110100010111: fc_kernel = 8'h11;
     14'b01110100011000: fc_kernel = 8'h04;
     14'b01110100011001: fc_kernel = 8'h00;
     14'b01110100011010: fc_kernel = 8'h02;
     14'b01110100011011: fc_kernel = 8'h01;
     14'b01110100011100: fc_kernel = 8'h00;
     14'b01110100011101: fc_kernel = 8'hf7;
     14'b01110100011110: fc_kernel = 8'hf7;
     14'b01110100011111: fc_kernel = 8'hfd;
     14'b01110100100000: fc_kernel = 8'h21;
     14'b01110100100001: fc_kernel = 8'h1a;
     14'b01110100100010: fc_kernel = 8'h0d;
     14'b01110100100011: fc_kernel = 8'h06;
     14'b01110100100100: fc_kernel = 8'h01;
     14'b01110100100101: fc_kernel = 8'h01;
     14'b01110100100110: fc_kernel = 8'hf7;
     14'b01110100100111: fc_kernel = 8'hf6;
     14'b01110100101000: fc_kernel = 8'h00;
     14'b01110100101001: fc_kernel = 8'hf0;
     14'b01110100101010: fc_kernel = 8'hd0;
     14'b01110100101011: fc_kernel = 8'hdc;
     14'b01110100101100: fc_kernel = 8'hf9;
     14'b01110100101101: fc_kernel = 8'h04;
     14'b01110100101110: fc_kernel = 8'h05;
     14'b01110100101111: fc_kernel = 8'h0d;
     14'b01110100110000: fc_kernel = 8'h0e;
     14'b01110100110001: fc_kernel = 8'h08;
     14'b01110100110010: fc_kernel = 8'h0d;
     14'b01110100110011: fc_kernel = 8'h06;
     14'b01110100110100: fc_kernel = 8'h06;
     14'b01110100110101: fc_kernel = 8'h00;
     14'b01110100110110: fc_kernel = 8'hfd;
     14'b01110100110111: fc_kernel = 8'hf5;
     14'b01110100111000: fc_kernel = 8'h1c;
     14'b01110100111001: fc_kernel = 8'h0c;
     14'b01110100111010: fc_kernel = 8'h05;
     14'b01110100111011: fc_kernel = 8'hfc;
     14'b01110100111100: fc_kernel = 8'hfc;
     14'b01110100111101: fc_kernel = 8'hfa;
     14'b01110100111110: fc_kernel = 8'hf5;
     14'b01110100111111: fc_kernel = 8'hfa;
     14'b01110101000000: fc_kernel = 8'hf8;
     14'b01110101000001: fc_kernel = 8'hea;
     14'b01110101000010: fc_kernel = 8'hdd;
     14'b01110101000011: fc_kernel = 8'he6;
     14'b01110101000100: fc_kernel = 8'hf5;
     14'b01110101000101: fc_kernel = 8'hfc;
     14'b01110101000110: fc_kernel = 8'h05;
     14'b01110101000111: fc_kernel = 8'h0e;
     14'b01110101001000: fc_kernel = 8'h0f;
     14'b01110101001001: fc_kernel = 8'h0e;
     14'b01110101001010: fc_kernel = 8'h10;
     14'b01110101001011: fc_kernel = 8'h07;
     14'b01110101001100: fc_kernel = 8'h03;
     14'b01110101001101: fc_kernel = 8'h02;
     14'b01110101001110: fc_kernel = 8'hf4;
     14'b01110101001111: fc_kernel = 8'hd5;
     14'b01110101010000: fc_kernel = 8'h09;
     14'b01110101010001: fc_kernel = 8'h00;
     14'b01110101010010: fc_kernel = 8'hfc;
     14'b01110101010011: fc_kernel = 8'hf9;
     14'b01110101010100: fc_kernel = 8'h01;
     14'b01110101010101: fc_kernel = 8'h02;
     14'b01110101010110: fc_kernel = 8'hfc;
     14'b01110101010111: fc_kernel = 8'hf7;
     14'b01110101011000: fc_kernel = 8'hee;
     14'b01110101011001: fc_kernel = 8'he3;
     14'b01110101011010: fc_kernel = 8'he6;
     14'b01110101011011: fc_kernel = 8'hf7;
     14'b01110101011100: fc_kernel = 8'hfb;
     14'b01110101011101: fc_kernel = 8'hfa;
     14'b01110101011110: fc_kernel = 8'h02;
     14'b01110101011111: fc_kernel = 8'h0d;
     14'b01110101100000: fc_kernel = 8'h0d;
     14'b01110101100001: fc_kernel = 8'h0c;
     14'b01110101100010: fc_kernel = 8'h09;
     14'b01110101100011: fc_kernel = 8'h04;
     14'b01110101100100: fc_kernel = 8'h02;
     14'b01110101100101: fc_kernel = 8'hf8;
     14'b01110101100110: fc_kernel = 8'hec;
     14'b01110101100111: fc_kernel = 8'hdc;
     14'b01110101101000: fc_kernel = 8'h00;
     14'b01110101101001: fc_kernel = 8'hfc;
     14'b01110101101010: fc_kernel = 8'hff;
     14'b01110101101011: fc_kernel = 8'hfd;
     14'b01110101101100: fc_kernel = 8'hf8;
     14'b01110101101101: fc_kernel = 8'hfb;
     14'b01110101101110: fc_kernel = 8'hfe;
     14'b01110101101111: fc_kernel = 8'hfb;
     14'b01110101110000: fc_kernel = 8'hec;
     14'b01110101110001: fc_kernel = 8'he9;
     14'b01110101110010: fc_kernel = 8'hf7;
     14'b01110101110011: fc_kernel = 8'hf8;
     14'b01110101110100: fc_kernel = 8'hfb;
     14'b01110101110101: fc_kernel = 8'h00;
     14'b01110101110110: fc_kernel = 8'h02;
     14'b01110101110111: fc_kernel = 8'h03;
     14'b01110101111000: fc_kernel = 8'h07;
     14'b01110101111001: fc_kernel = 8'h02;
     14'b01110101111010: fc_kernel = 8'h01;
     14'b01110101111011: fc_kernel = 8'hff;
     14'b01110101111100: fc_kernel = 8'hfb;
     14'b01110101111101: fc_kernel = 8'hf3;
     14'b01110101111110: fc_kernel = 8'hf2;
     14'b01110101111111: fc_kernel = 8'hf2;
     14'b01110110000000: fc_kernel = 8'h02;
     14'b01110110000001: fc_kernel = 8'h04;
     14'b01110110000010: fc_kernel = 8'h07;
     14'b01110110000011: fc_kernel = 8'h00;
     14'b01110110000100: fc_kernel = 8'hf4;
     14'b01110110000101: fc_kernel = 8'hf8;
     14'b01110110000110: fc_kernel = 8'hf5;
     14'b01110110000111: fc_kernel = 8'hef;
     14'b01110110001000: fc_kernel = 8'he9;
     14'b01110110001001: fc_kernel = 8'hf0;
     14'b01110110001010: fc_kernel = 8'hf2;
     14'b01110110001011: fc_kernel = 8'hfa;
     14'b01110110001100: fc_kernel = 8'h00;
     14'b01110110001101: fc_kernel = 8'hff;
     14'b01110110001110: fc_kernel = 8'h00;
     14'b01110110001111: fc_kernel = 8'h00;
     14'b01110110010000: fc_kernel = 8'hfe;
     14'b01110110010001: fc_kernel = 8'h00;
     14'b01110110010010: fc_kernel = 8'hfc;
     14'b01110110010011: fc_kernel = 8'hfe;
     14'b01110110010100: fc_kernel = 8'hf6;
     14'b01110110010101: fc_kernel = 8'hea;
     14'b01110110010110: fc_kernel = 8'hec;
     14'b01110110010111: fc_kernel = 8'hf3;
     14'b01110110011000: fc_kernel = 8'h06;
     14'b01110110011001: fc_kernel = 8'h00;
     14'b01110110011010: fc_kernel = 8'hff;
     14'b01110110011011: fc_kernel = 8'hfb;
     14'b01110110011100: fc_kernel = 8'hee;
     14'b01110110011101: fc_kernel = 8'hf0;
     14'b01110110011110: fc_kernel = 8'hee;
     14'b01110110011111: fc_kernel = 8'hec;
     14'b01110110100000: fc_kernel = 8'he6;
     14'b01110110100001: fc_kernel = 8'hec;
     14'b01110110100010: fc_kernel = 8'hf6;
     14'b01110110100011: fc_kernel = 8'h00;
     14'b01110110100100: fc_kernel = 8'h03;
     14'b01110110100101: fc_kernel = 8'hf8;
     14'b01110110100110: fc_kernel = 8'hf9;
     14'b01110110100111: fc_kernel = 8'hf2;
     14'b01110110101000: fc_kernel = 8'hf6;
     14'b01110110101001: fc_kernel = 8'hf7;
     14'b01110110101010: fc_kernel = 8'hf9;
     14'b01110110101011: fc_kernel = 8'hf9;
     14'b01110110101100: fc_kernel = 8'heb;
     14'b01110110101101: fc_kernel = 8'he8;
     14'b01110110101110: fc_kernel = 8'he5;
     14'b01110110101111: fc_kernel = 8'hf3;
     14'b01110110110000: fc_kernel = 8'h00;
     14'b01110110110001: fc_kernel = 8'hfd;
     14'b01110110110010: fc_kernel = 8'hf0;
     14'b01110110110011: fc_kernel = 8'hef;
     14'b01110110110100: fc_kernel = 8'hdc;
     14'b01110110110101: fc_kernel = 8'he6;
     14'b01110110110110: fc_kernel = 8'hee;
     14'b01110110110111: fc_kernel = 8'hed;
     14'b01110110111000: fc_kernel = 8'hea;
     14'b01110110111001: fc_kernel = 8'hed;
     14'b01110110111010: fc_kernel = 8'hf3;
     14'b01110110111011: fc_kernel = 8'hfe;
     14'b01110110111100: fc_kernel = 8'hfe;
     14'b01110110111101: fc_kernel = 8'hf8;
     14'b01110110111110: fc_kernel = 8'hec;
     14'b01110110111111: fc_kernel = 8'hec;
     14'b01110111000000: fc_kernel = 8'heb;
     14'b01110111000001: fc_kernel = 8'he5;
     14'b01110111000010: fc_kernel = 8'hee;
     14'b01110111000011: fc_kernel = 8'he6;
     14'b01110111000100: fc_kernel = 8'he1;
     14'b01110111000101: fc_kernel = 8'he1;
     14'b01110111000110: fc_kernel = 8'he9;
     14'b01110111000111: fc_kernel = 8'hf2;
     14'b01110111001000: fc_kernel = 8'hf1;
     14'b01110111001001: fc_kernel = 8'he2;
     14'b01110111001010: fc_kernel = 8'he4;
     14'b01110111001011: fc_kernel = 8'he5;
     14'b01110111001100: fc_kernel = 8'hdb;
     14'b01110111001101: fc_kernel = 8'he7;
     14'b01110111001110: fc_kernel = 8'hf3;
     14'b01110111001111: fc_kernel = 8'hf1;
     14'b01110111010000: fc_kernel = 8'hef;
     14'b01110111010001: fc_kernel = 8'hf7;
     14'b01110111010010: fc_kernel = 8'hfb;
     14'b01110111010011: fc_kernel = 8'hfd;
     14'b01110111010100: fc_kernel = 8'hfb;
     14'b01110111010101: fc_kernel = 8'hfc;
     14'b01110111010110: fc_kernel = 8'hf6;
     14'b01110111010111: fc_kernel = 8'heb;
     14'b01110111011000: fc_kernel = 8'hee;
     14'b01110111011001: fc_kernel = 8'hea;
     14'b01110111011010: fc_kernel = 8'he5;
     14'b01110111011011: fc_kernel = 8'he5;
     14'b01110111011100: fc_kernel = 8'he6;
     14'b01110111011101: fc_kernel = 8'hda;
     14'b01110111011110: fc_kernel = 8'he8;
     14'b01110111011111: fc_kernel = 8'hf6;
     14'b01110111100000: fc_kernel = 8'hda;
     14'b01110111100001: fc_kernel = 8'hdc;
     14'b01110111100010: fc_kernel = 8'he8;
     14'b01110111100011: fc_kernel = 8'hec;
     14'b01110111100100: fc_kernel = 8'hf1;
     14'b01110111100101: fc_kernel = 8'hf6;
     14'b01110111100110: fc_kernel = 8'hf4;
     14'b01110111100111: fc_kernel = 8'hf1;
     14'b01110111101000: fc_kernel = 8'hf1;
     14'b01110111101001: fc_kernel = 8'hf7;
     14'b01110111101010: fc_kernel = 8'hf7;
     14'b01110111101011: fc_kernel = 8'hf3;
     14'b01110111101100: fc_kernel = 8'hf4;
     14'b01110111101101: fc_kernel = 8'hf7;
     14'b01110111101110: fc_kernel = 8'hf7;
     14'b01110111101111: fc_kernel = 8'hee;
     14'b01110111110000: fc_kernel = 8'he8;
     14'b01110111110001: fc_kernel = 8'he9;
     14'b01110111110010: fc_kernel = 8'he9;
     14'b01110111110011: fc_kernel = 8'hdf;
     14'b01110111110100: fc_kernel = 8'hdd;
     14'b01110111110101: fc_kernel = 8'hcc;
     14'b01110111110110: fc_kernel = 8'hdd;
     14'b01110111110111: fc_kernel = 8'hfa;
     14'b01110111111000: fc_kernel = 8'hdb;
     14'b01110111111001: fc_kernel = 8'he1;
     14'b01110111111010: fc_kernel = 8'hf5;
     14'b01110111111011: fc_kernel = 8'h01;
     14'b01110111111100: fc_kernel = 8'h08;
     14'b01110111111101: fc_kernel = 8'h00;
     14'b01110111111110: fc_kernel = 8'hf4;
     14'b01110111111111: fc_kernel = 8'hf1;
     14'b01111000000000: fc_kernel = 8'hf1;
     14'b01111000000001: fc_kernel = 8'hf0;
     14'b01111000000010: fc_kernel = 8'hed;
     14'b01111000000011: fc_kernel = 8'hf2;
     14'b01111000000100: fc_kernel = 8'hf3;
     14'b01111000000101: fc_kernel = 8'hfa;
     14'b01111000000110: fc_kernel = 8'hf8;
     14'b01111000000111: fc_kernel = 8'hee;
     14'b01111000001000: fc_kernel = 8'he8;
     14'b01111000001001: fc_kernel = 8'he6;
     14'b01111000001010: fc_kernel = 8'hdf;
     14'b01111000001011: fc_kernel = 8'he0;
     14'b01111000001100: fc_kernel = 8'hd7;
     14'b01111000001101: fc_kernel = 8'hd4;
     14'b01111000001110: fc_kernel = 8'hca;
     14'b01111000001111: fc_kernel = 8'he5;
     14'b01111000010000: fc_kernel = 8'hea;
     14'b01111000010001: fc_kernel = 8'hfc;
     14'b01111000010010: fc_kernel = 8'h0d;
     14'b01111000010011: fc_kernel = 8'h12;
     14'b01111000010100: fc_kernel = 8'h0e;
     14'b01111000010101: fc_kernel = 8'h0b;
     14'b01111000010110: fc_kernel = 8'h00;
     14'b01111000010111: fc_kernel = 8'hfd;
     14'b01111000011000: fc_kernel = 8'hfc;
     14'b01111000011001: fc_kernel = 8'hfe;
     14'b01111000011010: fc_kernel = 8'hfe;
     14'b01111000011011: fc_kernel = 8'hfd;
     14'b01111000011100: fc_kernel = 8'hfe;
     14'b01111000011101: fc_kernel = 8'hf9;
     14'b01111000011110: fc_kernel = 8'hf6;
     14'b01111000011111: fc_kernel = 8'hf8;
     14'b01111000100000: fc_kernel = 8'hef;
     14'b01111000100001: fc_kernel = 8'hee;
     14'b01111000100010: fc_kernel = 8'he6;
     14'b01111000100011: fc_kernel = 8'he4;
     14'b01111000100100: fc_kernel = 8'he8;
     14'b01111000100101: fc_kernel = 8'hde;
     14'b01111000100110: fc_kernel = 8'hd0;
     14'b01111000100111: fc_kernel = 8'hdd;
     14'b01111000101000: fc_kernel = 8'hfa;
     14'b01111000101001: fc_kernel = 8'h0f;
     14'b01111000101010: fc_kernel = 8'h11;
     14'b01111000101011: fc_kernel = 8'h11;
     14'b01111000101100: fc_kernel = 8'h08;
     14'b01111000101101: fc_kernel = 8'h03;
     14'b01111000101110: fc_kernel = 8'h0c;
     14'b01111000101111: fc_kernel = 8'h0a;
     14'b01111000110000: fc_kernel = 8'h0d;
     14'b01111000110001: fc_kernel = 8'h0d;
     14'b01111000110010: fc_kernel = 8'h10;
     14'b01111000110011: fc_kernel = 8'h08;
     14'b01111000110100: fc_kernel = 8'h0d;
     14'b01111000110101: fc_kernel = 8'h0c;
     14'b01111000110110: fc_kernel = 8'h0c;
     14'b01111000110111: fc_kernel = 8'h09;
     14'b01111000111000: fc_kernel = 8'h0b;
     14'b01111000111001: fc_kernel = 8'h02;
     14'b01111000111010: fc_kernel = 8'hf7;
     14'b01111000111011: fc_kernel = 8'hf1;
     14'b01111000111100: fc_kernel = 8'hf8;
     14'b01111000111101: fc_kernel = 8'he9;
     14'b01111000111110: fc_kernel = 8'hdb;
     14'b01111000111111: fc_kernel = 8'hea;
     14'b10000000000000: fc_kernel = 8'he0;
     14'b10000000000001: fc_kernel = 8'hd9;
     14'b10000000000010: fc_kernel = 8'hee;
     14'b10000000000011: fc_kernel = 8'h0a;
     14'b10000000000100: fc_kernel = 8'h12;
     14'b10000000000101: fc_kernel = 8'hf2;
     14'b10000000000110: fc_kernel = 8'he5;
     14'b10000000000111: fc_kernel = 8'he0;
     14'b10000000001000: fc_kernel = 8'hde;
     14'b10000000001001: fc_kernel = 8'hda;
     14'b10000000001010: fc_kernel = 8'hc8;
     14'b10000000001011: fc_kernel = 8'hca;
     14'b10000000001100: fc_kernel = 8'he2;
     14'b10000000001101: fc_kernel = 8'hdc;
     14'b10000000001110: fc_kernel = 8'hd0;
     14'b10000000001111: fc_kernel = 8'he5;
     14'b10000000010000: fc_kernel = 8'hf5;
     14'b10000000010001: fc_kernel = 8'hde;
     14'b10000000010010: fc_kernel = 8'he0;
     14'b10000000010011: fc_kernel = 8'he0;
     14'b10000000010100: fc_kernel = 8'hf5;
     14'b10000000010101: fc_kernel = 8'hfb;
     14'b10000000010110: fc_kernel = 8'hf6;
     14'b10000000010111: fc_kernel = 8'hf6;
     14'b10000000011000: fc_kernel = 8'hed;
     14'b10000000011001: fc_kernel = 8'he0;
     14'b10000000011010: fc_kernel = 8'h03;
     14'b10000000011011: fc_kernel = 8'hf6;
     14'b10000000011100: fc_kernel = 8'hee;
     14'b10000000011101: fc_kernel = 8'he5;
     14'b10000000011110: fc_kernel = 8'he8;
     14'b10000000011111: fc_kernel = 8'hf2;
     14'b10000000100000: fc_kernel = 8'hf8;
     14'b10000000100001: fc_kernel = 8'hf0;
     14'b10000000100010: fc_kernel = 8'hfb;
     14'b10000000100011: fc_kernel = 8'hf4;
     14'b10000000100100: fc_kernel = 8'hf9;
     14'b10000000100101: fc_kernel = 8'hf1;
     14'b10000000100110: fc_kernel = 8'hee;
     14'b10000000100111: fc_kernel = 8'hfa;
     14'b10000000101000: fc_kernel = 8'hfc;
     14'b10000000101001: fc_kernel = 8'hf2;
     14'b10000000101010: fc_kernel = 8'hf6;
     14'b10000000101011: fc_kernel = 8'hfc;
     14'b10000000101100: fc_kernel = 8'h09;
     14'b10000000101101: fc_kernel = 8'h0c;
     14'b10000000101110: fc_kernel = 8'hff;
     14'b10000000101111: fc_kernel = 8'hf8;
     14'b10000000110000: fc_kernel = 8'hfa;
     14'b10000000110001: fc_kernel = 8'hf0;
     14'b10000000110010: fc_kernel = 8'he4;
     14'b10000000110011: fc_kernel = 8'hea;
     14'b10000000110100: fc_kernel = 8'hef;
     14'b10000000110101: fc_kernel = 8'hf8;
     14'b10000000110110: fc_kernel = 8'hfd;
     14'b10000000110111: fc_kernel = 8'hff;
     14'b10000000111000: fc_kernel = 8'hfe;
     14'b10000000111001: fc_kernel = 8'h03;
     14'b10000000111010: fc_kernel = 8'hfe;
     14'b10000000111011: fc_kernel = 8'h06;
     14'b10000000111100: fc_kernel = 8'h07;
     14'b10000000111101: fc_kernel = 8'h07;
     14'b10000000111110: fc_kernel = 8'h04;
     14'b10000000111111: fc_kernel = 8'h03;
     14'b10000001000000: fc_kernel = 8'h01;
     14'b10000001000001: fc_kernel = 8'h06;
     14'b10000001000010: fc_kernel = 8'h03;
     14'b10000001000011: fc_kernel = 8'h03;
     14'b10000001000100: fc_kernel = 8'h00;
     14'b10000001000101: fc_kernel = 8'h01;
     14'b10000001000110: fc_kernel = 8'h08;
     14'b10000001000111: fc_kernel = 8'h18;
     14'b10000001001000: fc_kernel = 8'h00;
     14'b10000001001001: fc_kernel = 8'he2;
     14'b10000001001010: fc_kernel = 8'hdf;
     14'b10000001001011: fc_kernel = 8'hdf;
     14'b10000001001100: fc_kernel = 8'hf5;
     14'b10000001001101: fc_kernel = 8'hff;
     14'b10000001001110: fc_kernel = 8'h03;
     14'b10000001001111: fc_kernel = 8'hf8;
     14'b10000001010000: fc_kernel = 8'hfc;
     14'b10000001010001: fc_kernel = 8'h01;
     14'b10000001010010: fc_kernel = 8'h08;
     14'b10000001010011: fc_kernel = 8'h07;
     14'b10000001010100: fc_kernel = 8'h08;
     14'b10000001010101: fc_kernel = 8'h07;
     14'b10000001010110: fc_kernel = 8'h03;
     14'b10000001010111: fc_kernel = 8'h06;
     14'b10000001011000: fc_kernel = 8'h01;
     14'b10000001011001: fc_kernel = 8'h02;
     14'b10000001011010: fc_kernel = 8'h03;
     14'b10000001011011: fc_kernel = 8'h02;
     14'b10000001011100: fc_kernel = 8'hf8;
     14'b10000001011101: fc_kernel = 8'hf5;
     14'b10000001011110: fc_kernel = 8'hfe;
     14'b10000001011111: fc_kernel = 8'h12;
     14'b10000001100000: fc_kernel = 8'hed;
     14'b10000001100001: fc_kernel = 8'hef;
     14'b10000001100010: fc_kernel = 8'heb;
     14'b10000001100011: fc_kernel = 8'hf0;
     14'b10000001100100: fc_kernel = 8'hf5;
     14'b10000001100101: fc_kernel = 8'hfd;
     14'b10000001100110: fc_kernel = 8'hff;
     14'b10000001100111: fc_kernel = 8'hf9;
     14'b10000001101000: fc_kernel = 8'hfd;
     14'b10000001101001: fc_kernel = 8'h01;
     14'b10000001101010: fc_kernel = 8'hff;
     14'b10000001101011: fc_kernel = 8'hfd;
     14'b10000001101100: fc_kernel = 8'h01;
     14'b10000001101101: fc_kernel = 8'h00;
     14'b10000001101110: fc_kernel = 8'h04;
     14'b10000001101111: fc_kernel = 8'h00;
     14'b10000001110000: fc_kernel = 8'h00;
     14'b10000001110001: fc_kernel = 8'h02;
     14'b10000001110010: fc_kernel = 8'h09;
     14'b10000001110011: fc_kernel = 8'hfd;
     14'b10000001110100: fc_kernel = 8'h00;
     14'b10000001110101: fc_kernel = 8'hfd;
     14'b10000001110110: fc_kernel = 8'h00;
     14'b10000001110111: fc_kernel = 8'h0c;
     14'b10000001111000: fc_kernel = 8'he7;
     14'b10000001111001: fc_kernel = 8'hf7;
     14'b10000001111010: fc_kernel = 8'hf9;
     14'b10000001111011: fc_kernel = 8'hf9;
     14'b10000001111100: fc_kernel = 8'hf9;
     14'b10000001111101: fc_kernel = 8'h01;
     14'b10000001111110: fc_kernel = 8'h00;
     14'b10000001111111: fc_kernel = 8'hfe;
     14'b10000010000000: fc_kernel = 8'hfd;
     14'b10000010000001: fc_kernel = 8'hfe;
     14'b10000010000010: fc_kernel = 8'h02;
     14'b10000010000011: fc_kernel = 8'h00;
     14'b10000010000100: fc_kernel = 8'h00;
     14'b10000010000101: fc_kernel = 8'h07;
     14'b10000010000110: fc_kernel = 8'h04;
     14'b10000010000111: fc_kernel = 8'hfd;
     14'b10000010001000: fc_kernel = 8'h00;
     14'b10000010001001: fc_kernel = 8'h01;
     14'b10000010001010: fc_kernel = 8'h03;
     14'b10000010001011: fc_kernel = 8'h01;
     14'b10000010001100: fc_kernel = 8'h01;
     14'b10000010001101: fc_kernel = 8'hfe;
     14'b10000010001110: fc_kernel = 8'h00;
     14'b10000010001111: fc_kernel = 8'h01;
     14'b10000010010000: fc_kernel = 8'h07;
     14'b10000010010001: fc_kernel = 8'hfc;
     14'b10000010010010: fc_kernel = 8'hfe;
     14'b10000010010011: fc_kernel = 8'hfb;
     14'b10000010010100: fc_kernel = 8'h01;
     14'b10000010010101: fc_kernel = 8'h03;
     14'b10000010010110: fc_kernel = 8'h02;
     14'b10000010010111: fc_kernel = 8'h06;
     14'b10000010011000: fc_kernel = 8'h00;
     14'b10000010011001: fc_kernel = 8'hff;
     14'b10000010011010: fc_kernel = 8'h02;
     14'b10000010011011: fc_kernel = 8'h02;
     14'b10000010011100: fc_kernel = 8'hfe;
     14'b10000010011101: fc_kernel = 8'hff;
     14'b10000010011110: fc_kernel = 8'h01;
     14'b10000010011111: fc_kernel = 8'h01;
     14'b10000010100000: fc_kernel = 8'h03;
     14'b10000010100001: fc_kernel = 8'h03;
     14'b10000010100010: fc_kernel = 8'h04;
     14'b10000010100011: fc_kernel = 8'h02;
     14'b10000010100100: fc_kernel = 8'h01;
     14'b10000010100101: fc_kernel = 8'h06;
     14'b10000010100110: fc_kernel = 8'h09;
     14'b10000010100111: fc_kernel = 8'h11;
     14'b10000010101000: fc_kernel = 8'hf9;
     14'b10000010101001: fc_kernel = 8'h01;
     14'b10000010101010: fc_kernel = 8'hfd;
     14'b10000010101011: fc_kernel = 8'h00;
     14'b10000010101100: fc_kernel = 8'h07;
     14'b10000010101101: fc_kernel = 8'h03;
     14'b10000010101110: fc_kernel = 8'h02;
     14'b10000010101111: fc_kernel = 8'h01;
     14'b10000010110000: fc_kernel = 8'h07;
     14'b10000010110001: fc_kernel = 8'h02;
     14'b10000010110010: fc_kernel = 8'h00;
     14'b10000010110011: fc_kernel = 8'hfa;
     14'b10000010110100: fc_kernel = 8'hf8;
     14'b10000010110101: fc_kernel = 8'hf7;
     14'b10000010110110: fc_kernel = 8'hfc;
     14'b10000010110111: fc_kernel = 8'hff;
     14'b10000010111000: fc_kernel = 8'h00;
     14'b10000010111001: fc_kernel = 8'h01;
     14'b10000010111010: fc_kernel = 8'h07;
     14'b10000010111011: fc_kernel = 8'h07;
     14'b10000010111100: fc_kernel = 8'h09;
     14'b10000010111101: fc_kernel = 8'h04;
     14'b10000010111110: fc_kernel = 8'h09;
     14'b10000010111111: fc_kernel = 8'h09;
     14'b10000011000000: fc_kernel = 8'he8;
     14'b10000011000001: fc_kernel = 8'hfc;
     14'b10000011000010: fc_kernel = 8'hfa;
     14'b10000011000011: fc_kernel = 8'h05;
     14'b10000011000100: fc_kernel = 8'h00;
     14'b10000011000101: fc_kernel = 8'h05;
     14'b10000011000110: fc_kernel = 8'h07;
     14'b10000011000111: fc_kernel = 8'h06;
     14'b10000011001000: fc_kernel = 8'h07;
     14'b10000011001001: fc_kernel = 8'h09;
     14'b10000011001010: fc_kernel = 8'h0e;
     14'b10000011001011: fc_kernel = 8'h08;
     14'b10000011001100: fc_kernel = 8'hfa;
     14'b10000011001101: fc_kernel = 8'hec;
     14'b10000011001110: fc_kernel = 8'hf3;
     14'b10000011001111: fc_kernel = 8'h00;
     14'b10000011010000: fc_kernel = 8'h02;
     14'b10000011010001: fc_kernel = 8'h03;
     14'b10000011010010: fc_kernel = 8'h02;
     14'b10000011010011: fc_kernel = 8'h01;
     14'b10000011010100: fc_kernel = 8'h02;
     14'b10000011010101: fc_kernel = 8'h01;
     14'b10000011010110: fc_kernel = 8'hfa;
     14'b10000011010111: fc_kernel = 8'hf0;
     14'b10000011011000: fc_kernel = 8'he8;
     14'b10000011011001: fc_kernel = 8'hf8;
     14'b10000011011010: fc_kernel = 8'hfc;
     14'b10000011011011: fc_kernel = 8'h01;
     14'b10000011011100: fc_kernel = 8'h05;
     14'b10000011011101: fc_kernel = 8'h08;
     14'b10000011011110: fc_kernel = 8'h09;
     14'b10000011011111: fc_kernel = 8'h0a;
     14'b10000011100000: fc_kernel = 8'h07;
     14'b10000011100001: fc_kernel = 8'h09;
     14'b10000011100010: fc_kernel = 8'h05;
     14'b10000011100011: fc_kernel = 8'h07;
     14'b10000011100100: fc_kernel = 8'h01;
     14'b10000011100101: fc_kernel = 8'hf8;
     14'b10000011100110: fc_kernel = 8'hf4;
     14'b10000011100111: fc_kernel = 8'hf8;
     14'b10000011101000: fc_kernel = 8'h00;
     14'b10000011101001: fc_kernel = 8'h07;
     14'b10000011101010: fc_kernel = 8'h06;
     14'b10000011101011: fc_kernel = 8'h08;
     14'b10000011101100: fc_kernel = 8'h06;
     14'b10000011101101: fc_kernel = 8'h08;
     14'b10000011101110: fc_kernel = 8'h01;
     14'b10000011101111: fc_kernel = 8'hf0;
     14'b10000011110000: fc_kernel = 8'hff;
     14'b10000011110001: fc_kernel = 8'h00;
     14'b10000011110010: fc_kernel = 8'h05;
     14'b10000011110011: fc_kernel = 8'h04;
     14'b10000011110100: fc_kernel = 8'h08;
     14'b10000011110101: fc_kernel = 8'h04;
     14'b10000011110110: fc_kernel = 8'h0a;
     14'b10000011110111: fc_kernel = 8'h08;
     14'b10000011111000: fc_kernel = 8'h00;
     14'b10000011111001: fc_kernel = 8'hff;
     14'b10000011111010: fc_kernel = 8'hfe;
     14'b10000011111011: fc_kernel = 8'h05;
     14'b10000011111100: fc_kernel = 8'h06;
     14'b10000011111101: fc_kernel = 8'hfe;
     14'b10000011111110: fc_kernel = 8'hf9;
     14'b10000011111111: fc_kernel = 8'hfb;
     14'b10000100000000: fc_kernel = 8'hfe;
     14'b10000100000001: fc_kernel = 8'h03;
     14'b10000100000010: fc_kernel = 8'h04;
     14'b10000100000011: fc_kernel = 8'h0e;
     14'b10000100000100: fc_kernel = 8'h0f;
     14'b10000100000101: fc_kernel = 8'h12;
     14'b10000100000110: fc_kernel = 8'h10;
     14'b10000100000111: fc_kernel = 8'h04;
     14'b10000100001000: fc_kernel = 8'h03;
     14'b10000100001001: fc_kernel = 8'h00;
     14'b10000100001010: fc_kernel = 8'h06;
     14'b10000100001011: fc_kernel = 8'h05;
     14'b10000100001100: fc_kernel = 8'h03;
     14'b10000100001101: fc_kernel = 8'h06;
     14'b10000100001110: fc_kernel = 8'h00;
     14'b10000100001111: fc_kernel = 8'h00;
     14'b10000100010000: fc_kernel = 8'hf9;
     14'b10000100010001: fc_kernel = 8'h00;
     14'b10000100010010: fc_kernel = 8'h07;
     14'b10000100010011: fc_kernel = 8'h09;
     14'b10000100010100: fc_kernel = 8'h07;
     14'b10000100010101: fc_kernel = 8'h00;
     14'b10000100010110: fc_kernel = 8'hfe;
     14'b10000100010111: fc_kernel = 8'h01;
     14'b10000100011000: fc_kernel = 8'hfc;
     14'b10000100011001: fc_kernel = 8'h02;
     14'b10000100011010: fc_kernel = 8'h00;
     14'b10000100011011: fc_kernel = 8'h01;
     14'b10000100011100: fc_kernel = 8'h03;
     14'b10000100011101: fc_kernel = 8'h0f;
     14'b10000100011110: fc_kernel = 8'h14;
     14'b10000100011111: fc_kernel = 8'h03;
     14'b10000100100000: fc_kernel = 8'hfc;
     14'b10000100100001: fc_kernel = 8'hf6;
     14'b10000100100010: fc_kernel = 8'hfc;
     14'b10000100100011: fc_kernel = 8'hff;
     14'b10000100100100: fc_kernel = 8'hfd;
     14'b10000100100101: fc_kernel = 8'hf3;
     14'b10000100100110: fc_kernel = 8'hf7;
     14'b10000100100111: fc_kernel = 8'hf8;
     14'b10000100101000: fc_kernel = 8'hf8;
     14'b10000100101001: fc_kernel = 8'h03;
     14'b10000100101010: fc_kernel = 8'h08;
     14'b10000100101011: fc_kernel = 8'h08;
     14'b10000100101100: fc_kernel = 8'h05;
     14'b10000100101101: fc_kernel = 8'h00;
     14'b10000100101110: fc_kernel = 8'hfc;
     14'b10000100101111: fc_kernel = 8'hfa;
     14'b10000100110000: fc_kernel = 8'hfa;
     14'b10000100110001: fc_kernel = 8'hfe;
     14'b10000100110010: fc_kernel = 8'hfd;
     14'b10000100110011: fc_kernel = 8'hfc;
     14'b10000100110100: fc_kernel = 8'hf7;
     14'b10000100110101: fc_kernel = 8'hf9;
     14'b10000100110110: fc_kernel = 8'hfc;
     14'b10000100110111: fc_kernel = 8'h00;
     14'b10000100111000: fc_kernel = 8'hfc;
     14'b10000100111001: fc_kernel = 8'he2;
     14'b10000100111010: fc_kernel = 8'heb;
     14'b10000100111011: fc_kernel = 8'hf6;
     14'b10000100111100: fc_kernel = 8'hf4;
     14'b10000100111101: fc_kernel = 8'hef;
     14'b10000100111110: fc_kernel = 8'hf1;
     14'b10000100111111: fc_kernel = 8'hf4;
     14'b10000101000000: fc_kernel = 8'hff;
     14'b10000101000001: fc_kernel = 8'h01;
     14'b10000101000010: fc_kernel = 8'h0c;
     14'b10000101000011: fc_kernel = 8'h07;
     14'b10000101000100: fc_kernel = 8'h07;
     14'b10000101000101: fc_kernel = 8'h02;
     14'b10000101000110: fc_kernel = 8'hfc;
     14'b10000101000111: fc_kernel = 8'hf9;
     14'b10000101001000: fc_kernel = 8'hfc;
     14'b10000101001001: fc_kernel = 8'hff;
     14'b10000101001010: fc_kernel = 8'hf2;
     14'b10000101001011: fc_kernel = 8'hf7;
     14'b10000101001100: fc_kernel = 8'hf0;
     14'b10000101001101: fc_kernel = 8'heb;
     14'b10000101001110: fc_kernel = 8'he7;
     14'b10000101001111: fc_kernel = 8'hf5;
     14'b10000101010000: fc_kernel = 8'hf3;
     14'b10000101010001: fc_kernel = 8'hf7;
     14'b10000101010010: fc_kernel = 8'hde;
     14'b10000101010011: fc_kernel = 8'he7;
     14'b10000101010100: fc_kernel = 8'hf5;
     14'b10000101010101: fc_kernel = 8'hf7;
     14'b10000101010110: fc_kernel = 8'hfb;
     14'b10000101010111: fc_kernel = 8'h00;
     14'b10000101011000: fc_kernel = 8'hf8;
     14'b10000101011001: fc_kernel = 8'h00;
     14'b10000101011010: fc_kernel = 8'h04;
     14'b10000101011011: fc_kernel = 8'h07;
     14'b10000101011100: fc_kernel = 8'h02;
     14'b10000101011101: fc_kernel = 8'hff;
     14'b10000101011110: fc_kernel = 8'hfc;
     14'b10000101011111: fc_kernel = 8'hfa;
     14'b10000101100000: fc_kernel = 8'hf9;
     14'b10000101100001: fc_kernel = 8'hf5;
     14'b10000101100010: fc_kernel = 8'hf6;
     14'b10000101100011: fc_kernel = 8'hed;
     14'b10000101100100: fc_kernel = 8'hf2;
     14'b10000101100101: fc_kernel = 8'hef;
     14'b10000101100110: fc_kernel = 8'hf4;
     14'b10000101100111: fc_kernel = 8'he9;
     14'b10000101101000: fc_kernel = 8'hf0;
     14'b10000101101001: fc_kernel = 8'hf0;
     14'b10000101101010: fc_kernel = 8'hd6;
     14'b10000101101011: fc_kernel = 8'he1;
     14'b10000101101100: fc_kernel = 8'hf4;
     14'b10000101101101: fc_kernel = 8'hfc;
     14'b10000101101110: fc_kernel = 8'h02;
     14'b10000101101111: fc_kernel = 8'h02;
     14'b10000101110000: fc_kernel = 8'h03;
     14'b10000101110001: fc_kernel = 8'h0c;
     14'b10000101110010: fc_kernel = 8'h0d;
     14'b10000101110011: fc_kernel = 8'h09;
     14'b10000101110100: fc_kernel = 8'hfc;
     14'b10000101110101: fc_kernel = 8'h00;
     14'b10000101110110: fc_kernel = 8'hfd;
     14'b10000101110111: fc_kernel = 8'h00;
     14'b10000101111000: fc_kernel = 8'hf6;
     14'b10000101111001: fc_kernel = 8'hf4;
     14'b10000101111010: fc_kernel = 8'hf4;
     14'b10000101111011: fc_kernel = 8'hf3;
     14'b10000101111100: fc_kernel = 8'hed;
     14'b10000101111101: fc_kernel = 8'hfa;
     14'b10000101111110: fc_kernel = 8'hf6;
     14'b10000101111111: fc_kernel = 8'hea;
     14'b10000110000000: fc_kernel = 8'hde;
     14'b10000110000001: fc_kernel = 8'hce;
     14'b10000110000010: fc_kernel = 8'he9;
     14'b10000110000011: fc_kernel = 8'hfb;
     14'b10000110000100: fc_kernel = 8'hf4;
     14'b10000110000101: fc_kernel = 8'hfc;
     14'b10000110000110: fc_kernel = 8'h01;
     14'b10000110000111: fc_kernel = 8'h01;
     14'b10000110001000: fc_kernel = 8'h07;
     14'b10000110001001: fc_kernel = 8'h07;
     14'b10000110001010: fc_kernel = 8'h07;
     14'b10000110001011: fc_kernel = 8'h06;
     14'b10000110001100: fc_kernel = 8'hf8;
     14'b10000110001101: fc_kernel = 8'hfc;
     14'b10000110001110: fc_kernel = 8'hfa;
     14'b10000110001111: fc_kernel = 8'hf7;
     14'b10000110010000: fc_kernel = 8'hf8;
     14'b10000110010001: fc_kernel = 8'hf9;
     14'b10000110010010: fc_kernel = 8'hf6;
     14'b10000110010011: fc_kernel = 8'hf3;
     14'b10000110010100: fc_kernel = 8'hf5;
     14'b10000110010101: fc_kernel = 8'hfe;
     14'b10000110010110: fc_kernel = 8'hfd;
     14'b10000110010111: fc_kernel = 8'heb;
     14'b10000110011000: fc_kernel = 8'hca;
     14'b10000110011001: fc_kernel = 8'hd6;
     14'b10000110011010: fc_kernel = 8'hf2;
     14'b10000110011011: fc_kernel = 8'hfe;
     14'b10000110011100: fc_kernel = 8'hfd;
     14'b10000110011101: fc_kernel = 8'hf9;
     14'b10000110011110: fc_kernel = 8'h00;
     14'b10000110011111: fc_kernel = 8'h01;
     14'b10000110100000: fc_kernel = 8'h05;
     14'b10000110100001: fc_kernel = 8'h07;
     14'b10000110100010: fc_kernel = 8'h03;
     14'b10000110100011: fc_kernel = 8'hfc;
     14'b10000110100100: fc_kernel = 8'hf3;
     14'b10000110100101: fc_kernel = 8'hf9;
     14'b10000110100110: fc_kernel = 8'hfb;
     14'b10000110100111: fc_kernel = 8'hfb;
     14'b10000110101000: fc_kernel = 8'hf8;
     14'b10000110101001: fc_kernel = 8'h00;
     14'b10000110101010: fc_kernel = 8'hfb;
     14'b10000110101011: fc_kernel = 8'hfd;
     14'b10000110101100: fc_kernel = 8'h02;
     14'b10000110101101: fc_kernel = 8'h08;
     14'b10000110101110: fc_kernel = 8'hfc;
     14'b10000110101111: fc_kernel = 8'he8;
     14'b10000110110000: fc_kernel = 8'hc0;
     14'b10000110110001: fc_kernel = 8'he1;
     14'b10000110110010: fc_kernel = 8'hf4;
     14'b10000110110011: fc_kernel = 8'hf8;
     14'b10000110110100: fc_kernel = 8'h00;
     14'b10000110110101: fc_kernel = 8'h03;
     14'b10000110110110: fc_kernel = 8'h03;
     14'b10000110110111: fc_kernel = 8'h03;
     14'b10000110111000: fc_kernel = 8'h02;
     14'b10000110111001: fc_kernel = 8'hfc;
     14'b10000110111010: fc_kernel = 8'hfc;
     14'b10000110111011: fc_kernel = 8'hff;
     14'b10000110111100: fc_kernel = 8'hfb;
     14'b10000110111101: fc_kernel = 8'hf7;
     14'b10000110111110: fc_kernel = 8'hf8;
     14'b10000110111111: fc_kernel = 8'hfa;
     14'b10000111000000: fc_kernel = 8'hff;
     14'b10000111000001: fc_kernel = 8'h02;
     14'b10000111000010: fc_kernel = 8'h01;
     14'b10000111000011: fc_kernel = 8'h01;
     14'b10000111000100: fc_kernel = 8'h00;
     14'b10000111000101: fc_kernel = 8'h09;
     14'b10000111000110: fc_kernel = 8'hfc;
     14'b10000111000111: fc_kernel = 8'hdf;
     14'b10000111001000: fc_kernel = 8'hd1;
     14'b10000111001001: fc_kernel = 8'he9;
     14'b10000111001010: fc_kernel = 8'hf3;
     14'b10000111001011: fc_kernel = 8'hfe;
     14'b10000111001100: fc_kernel = 8'h00;
     14'b10000111001101: fc_kernel = 8'h05;
     14'b10000111001110: fc_kernel = 8'h02;
     14'b10000111001111: fc_kernel = 8'h04;
     14'b10000111010000: fc_kernel = 8'h00;
     14'b10000111010001: fc_kernel = 8'h03;
     14'b10000111010010: fc_kernel = 8'h00;
     14'b10000111010011: fc_kernel = 8'hff;
     14'b10000111010100: fc_kernel = 8'h01;
     14'b10000111010101: fc_kernel = 8'hfe;
     14'b10000111010110: fc_kernel = 8'hfb;
     14'b10000111010111: fc_kernel = 8'hfa;
     14'b10000111011000: fc_kernel = 8'hf9;
     14'b10000111011001: fc_kernel = 8'hfc;
     14'b10000111011010: fc_kernel = 8'h01;
     14'b10000111011011: fc_kernel = 8'h01;
     14'b10000111011100: fc_kernel = 8'hff;
     14'b10000111011101: fc_kernel = 8'h02;
     14'b10000111011110: fc_kernel = 8'hf5;
     14'b10000111011111: fc_kernel = 8'hdd;
     14'b10000111100000: fc_kernel = 8'hd2;
     14'b10000111100001: fc_kernel = 8'hf5;
     14'b10000111100010: fc_kernel = 8'hfb;
     14'b10000111100011: fc_kernel = 8'hfc;
     14'b10000111100100: fc_kernel = 8'h06;
     14'b10000111100101: fc_kernel = 8'h04;
     14'b10000111100110: fc_kernel = 8'h00;
     14'b10000111100111: fc_kernel = 8'hfe;
     14'b10000111101000: fc_kernel = 8'h00;
     14'b10000111101001: fc_kernel = 8'hfe;
     14'b10000111101010: fc_kernel = 8'h00;
     14'b10000111101011: fc_kernel = 8'h06;
     14'b10000111101100: fc_kernel = 8'h02;
     14'b10000111101101: fc_kernel = 8'hfe;
     14'b10000111101110: fc_kernel = 8'h03;
     14'b10000111101111: fc_kernel = 8'h00;
     14'b10000111110000: fc_kernel = 8'h02;
     14'b10000111110001: fc_kernel = 8'hfe;
     14'b10000111110010: fc_kernel = 8'hff;
     14'b10000111110011: fc_kernel = 8'h01;
     14'b10000111110100: fc_kernel = 8'h03;
     14'b10000111110101: fc_kernel = 8'h09;
     14'b10000111110110: fc_kernel = 8'hf8;
     14'b10000111110111: fc_kernel = 8'he8;
     14'b10000111111000: fc_kernel = 8'hd8;
     14'b10000111111001: fc_kernel = 8'hf6;
     14'b10000111111010: fc_kernel = 8'hfa;
     14'b10000111111011: fc_kernel = 8'hf8;
     14'b10000111111100: fc_kernel = 8'hf9;
     14'b10000111111101: fc_kernel = 8'hfb;
     14'b10000111111110: fc_kernel = 8'h05;
     14'b10000111111111: fc_kernel = 8'h01;
     14'b10001000000000: fc_kernel = 8'h01;
     14'b10001000000001: fc_kernel = 8'h05;
     14'b10001000000010: fc_kernel = 8'h04;
     14'b10001000000011: fc_kernel = 8'h09;
     14'b10001000000100: fc_kernel = 8'h09;
     14'b10001000000101: fc_kernel = 8'h03;
     14'b10001000000110: fc_kernel = 8'h02;
     14'b10001000000111: fc_kernel = 8'h00;
     14'b10001000001000: fc_kernel = 8'h07;
     14'b10001000001001: fc_kernel = 8'h01;
     14'b10001000001010: fc_kernel = 8'h02;
     14'b10001000001011: fc_kernel = 8'h03;
     14'b10001000001100: fc_kernel = 8'h08;
     14'b10001000001101: fc_kernel = 8'hff;
     14'b10001000001110: fc_kernel = 8'h03;
     14'b10001000001111: fc_kernel = 8'he9;
     14'b10001000010000: fc_kernel = 8'hea;
     14'b10001000010001: fc_kernel = 8'heb;
     14'b10001000010010: fc_kernel = 8'hec;
     14'b10001000010011: fc_kernel = 8'hec;
     14'b10001000010100: fc_kernel = 8'hea;
     14'b10001000010101: fc_kernel = 8'hfb;
     14'b10001000010110: fc_kernel = 8'h01;
     14'b10001000010111: fc_kernel = 8'h02;
     14'b10001000011000: fc_kernel = 8'h02;
     14'b10001000011001: fc_kernel = 8'h04;
     14'b10001000011010: fc_kernel = 8'h0b;
     14'b10001000011011: fc_kernel = 8'h06;
     14'b10001000011100: fc_kernel = 8'h06;
     14'b10001000011101: fc_kernel = 8'h09;
     14'b10001000011110: fc_kernel = 8'h0a;
     14'b10001000011111: fc_kernel = 8'h07;
     14'b10001000100000: fc_kernel = 8'h03;
     14'b10001000100001: fc_kernel = 8'h0e;
     14'b10001000100010: fc_kernel = 8'h0b;
     14'b10001000100011: fc_kernel = 8'h01;
     14'b10001000100100: fc_kernel = 8'h00;
     14'b10001000100101: fc_kernel = 8'hfe;
     14'b10001000100110: fc_kernel = 8'hf5;
     14'b10001000100111: fc_kernel = 8'hda;
     14'b10001000101000: fc_kernel = 8'hee;
     14'b10001000101001: fc_kernel = 8'he2;
     14'b10001000101010: fc_kernel = 8'hd6;
     14'b10001000101011: fc_kernel = 8'hdc;
     14'b10001000101100: fc_kernel = 8'he4;
     14'b10001000101101: fc_kernel = 8'hf4;
     14'b10001000101110: fc_kernel = 8'hf6;
     14'b10001000101111: fc_kernel = 8'hf5;
     14'b10001000110000: fc_kernel = 8'hf7;
     14'b10001000110001: fc_kernel = 8'h00;
     14'b10001000110010: fc_kernel = 8'hfc;
     14'b10001000110011: fc_kernel = 8'hf7;
     14'b10001000110100: fc_kernel = 8'hfe;
     14'b10001000110101: fc_kernel = 8'h02;
     14'b10001000110110: fc_kernel = 8'h06;
     14'b10001000110111: fc_kernel = 8'hff;
     14'b10001000111000: fc_kernel = 8'h00;
     14'b10001000111001: fc_kernel = 8'h0a;
     14'b10001000111010: fc_kernel = 8'h05;
     14'b10001000111011: fc_kernel = 8'hf7;
     14'b10001000111100: fc_kernel = 8'hf2;
     14'b10001000111101: fc_kernel = 8'he9;
     14'b10001000111110: fc_kernel = 8'he1;
     14'b10001000111111: fc_kernel = 8'hd9;
     14'b10010000000000: fc_kernel = 8'hf1;
     14'b10010000000001: fc_kernel = 8'hf2;
     14'b10010000000010: fc_kernel = 8'heb;
     14'b10010000000011: fc_kernel = 8'he8;
     14'b10010000000100: fc_kernel = 8'he3;
     14'b10010000000101: fc_kernel = 8'hdf;
     14'b10010000000110: fc_kernel = 8'hfe;
     14'b10010000000111: fc_kernel = 8'he2;
     14'b10010000001000: fc_kernel = 8'hc8;
     14'b10010000001001: fc_kernel = 8'hbd;
     14'b10010000001010: fc_kernel = 8'had;
     14'b10010000001011: fc_kernel = 8'ha3;
     14'b10010000001100: fc_kernel = 8'h9b;
     14'b10010000001101: fc_kernel = 8'hbf;
     14'b10010000001110: fc_kernel = 8'hcc;
     14'b10010000001111: fc_kernel = 8'he1;
     14'b10010000010000: fc_kernel = 8'hee;
     14'b10010000010001: fc_kernel = 8'hf5;
     14'b10010000010010: fc_kernel = 8'hf2;
     14'b10010000010011: fc_kernel = 8'hf6;
     14'b10010000010100: fc_kernel = 8'hea;
     14'b10010000010101: fc_kernel = 8'heb;
     14'b10010000010110: fc_kernel = 8'hf1;
     14'b10010000010111: fc_kernel = 8'hf2;
     14'b10010000011000: fc_kernel = 8'hec;
     14'b10010000011001: fc_kernel = 8'he7;
     14'b10010000011010: fc_kernel = 8'he2;
     14'b10010000011011: fc_kernel = 8'hfa;
     14'b10010000011100: fc_kernel = 8'heb;
     14'b10010000011101: fc_kernel = 8'heb;
     14'b10010000011110: fc_kernel = 8'he5;
     14'b10010000011111: fc_kernel = 8'heb;
     14'b10010000100000: fc_kernel = 8'ha6;
     14'b10010000100001: fc_kernel = 8'ha0;
     14'b10010000100010: fc_kernel = 8'h87;
     14'b10010000100011: fc_kernel = 8'h98;
     14'b10010000100100: fc_kernel = 8'h94;
     14'b10010000100101: fc_kernel = 8'ha6;
     14'b10010000100110: fc_kernel = 8'hac;
     14'b10010000100111: fc_kernel = 8'hc6;
     14'b10010000101000: fc_kernel = 8'hd7;
     14'b10010000101001: fc_kernel = 8'hdf;
     14'b10010000101010: fc_kernel = 8'hd2;
     14'b10010000101011: fc_kernel = 8'hd2;
     14'b10010000101100: fc_kernel = 8'hdc;
     14'b10010000101101: fc_kernel = 8'hdf;
     14'b10010000101110: fc_kernel = 8'he0;
     14'b10010000101111: fc_kernel = 8'he9;
     14'b10010000110000: fc_kernel = 8'hdf;
     14'b10010000110001: fc_kernel = 8'hd3;
     14'b10010000110010: fc_kernel = 8'h08;
     14'b10010000110011: fc_kernel = 8'hdc;
     14'b10010000110100: fc_kernel = 8'he9;
     14'b10010000110101: fc_kernel = 8'hdc;
     14'b10010000110110: fc_kernel = 8'hb7;
     14'b10010000110111: fc_kernel = 8'haf;
     14'b10010000111000: fc_kernel = 8'hb9;
     14'b10010000111001: fc_kernel = 8'hdd;
     14'b10010000111010: fc_kernel = 8'he6;
     14'b10010000111011: fc_kernel = 8'heb;
     14'b10010000111100: fc_kernel = 8'he8;
     14'b10010000111101: fc_kernel = 8'hdf;
     14'b10010000111110: fc_kernel = 8'hde;
     14'b10010000111111: fc_kernel = 8'he1;
     14'b10010001000000: fc_kernel = 8'he3;
     14'b10010001000001: fc_kernel = 8'hdc;
     14'b10010001000010: fc_kernel = 8'hd2;
     14'b10010001000011: fc_kernel = 8'hc9;
     14'b10010001000100: fc_kernel = 8'hc1;
     14'b10010001000101: fc_kernel = 8'hce;
     14'b10010001000110: fc_kernel = 8'hd9;
     14'b10010001000111: fc_kernel = 8'he0;
     14'b10010001001000: fc_kernel = 8'hdc;
     14'b10010001001001: fc_kernel = 8'he3;
     14'b10010001001010: fc_kernel = 8'hfa;
     14'b10010001001011: fc_kernel = 8'hd1;
     14'b10010001001100: fc_kernel = 8'hcd;
     14'b10010001001101: fc_kernel = 8'hc1;
     14'b10010001001110: fc_kernel = 8'hd0;
     14'b10010001001111: fc_kernel = 8'he2;
     14'b10010001010000: fc_kernel = 8'hf6;
     14'b10010001010001: fc_kernel = 8'h00;
     14'b10010001010010: fc_kernel = 8'h04;
     14'b10010001010011: fc_kernel = 8'h07;
     14'b10010001010100: fc_kernel = 8'h0a;
     14'b10010001010101: fc_kernel = 8'h00;
     14'b10010001010110: fc_kernel = 8'hf7;
     14'b10010001010111: fc_kernel = 8'hfa;
     14'b10010001011000: fc_kernel = 8'hf7;
     14'b10010001011001: fc_kernel = 8'hf9;
     14'b10010001011010: fc_kernel = 8'hfa;
     14'b10010001011011: fc_kernel = 8'hf1;
     14'b10010001011100: fc_kernel = 8'hd3;
     14'b10010001011101: fc_kernel = 8'hb4;
     14'b10010001011110: fc_kernel = 8'hc5;
     14'b10010001011111: fc_kernel = 8'hd7;
     14'b10010001100000: fc_kernel = 8'hef;
     14'b10010001100001: fc_kernel = 8'hf3;
     14'b10010001100010: fc_kernel = 8'hcf;
     14'b10010001100011: fc_kernel = 8'hb2;
     14'b10010001100100: fc_kernel = 8'hd3;
     14'b10010001100101: fc_kernel = 8'he3;
     14'b10010001100110: fc_kernel = 8'hef;
     14'b10010001100111: fc_kernel = 8'hf6;
     14'b10010001101000: fc_kernel = 8'hff;
     14'b10010001101001: fc_kernel = 8'h09;
     14'b10010001101010: fc_kernel = 8'h12;
     14'b10010001101011: fc_kernel = 8'h0a;
     14'b10010001101100: fc_kernel = 8'h0c;
     14'b10010001101101: fc_kernel = 8'h0a;
     14'b10010001101110: fc_kernel = 8'h0b;
     14'b10010001101111: fc_kernel = 8'h06;
     14'b10010001110000: fc_kernel = 8'h0b;
     14'b10010001110001: fc_kernel = 8'h06;
     14'b10010001110010: fc_kernel = 8'h00;
     14'b10010001110011: fc_kernel = 8'hfd;
     14'b10010001110100: fc_kernel = 8'hef;
     14'b10010001110101: fc_kernel = 8'hdd;
     14'b10010001110110: fc_kernel = 8'hdc;
     14'b10010001110111: fc_kernel = 8'heb;
     14'b10010001111000: fc_kernel = 8'hdf;
     14'b10010001111001: fc_kernel = 8'hf7;
     14'b10010001111010: fc_kernel = 8'hc9;
     14'b10010001111011: fc_kernel = 8'hd7;
     14'b10010001111100: fc_kernel = 8'he6;
     14'b10010001111101: fc_kernel = 8'hed;
     14'b10010001111110: fc_kernel = 8'hf9;
     14'b10010001111111: fc_kernel = 8'hfa;
     14'b10010010000000: fc_kernel = 8'hfd;
     14'b10010010000001: fc_kernel = 8'hfe;
     14'b10010010000010: fc_kernel = 8'h03;
     14'b10010010000011: fc_kernel = 8'h0e;
     14'b10010010000100: fc_kernel = 8'h0d;
     14'b10010010000101: fc_kernel = 8'h08;
     14'b10010010000110: fc_kernel = 8'h0b;
     14'b10010010000111: fc_kernel = 8'h06;
     14'b10010010001000: fc_kernel = 8'h00;
     14'b10010010001001: fc_kernel = 8'h00;
     14'b10010010001010: fc_kernel = 8'h03;
     14'b10010010001011: fc_kernel = 8'hfd;
     14'b10010010001100: fc_kernel = 8'hf9;
     14'b10010010001101: fc_kernel = 8'hed;
     14'b10010010001110: fc_kernel = 8'he9;
     14'b10010010001111: fc_kernel = 8'he1;
     14'b10010010010000: fc_kernel = 8'hd4;
     14'b10010010010001: fc_kernel = 8'hdc;
     14'b10010010010010: fc_kernel = 8'he0;
     14'b10010010010011: fc_kernel = 8'hf0;
     14'b10010010010100: fc_kernel = 8'hf5;
     14'b10010010010101: fc_kernel = 8'hf7;
     14'b10010010010110: fc_kernel = 8'hfb;
     14'b10010010010111: fc_kernel = 8'hfc;
     14'b10010010011000: fc_kernel = 8'hff;
     14'b10010010011001: fc_kernel = 8'hfd;
     14'b10010010011010: fc_kernel = 8'h00;
     14'b10010010011011: fc_kernel = 8'h06;
     14'b10010010011100: fc_kernel = 8'h12;
     14'b10010010011101: fc_kernel = 8'h0c;
     14'b10010010011110: fc_kernel = 8'h0c;
     14'b10010010011111: fc_kernel = 8'h05;
     14'b10010010100000: fc_kernel = 8'h06;
     14'b10010010100001: fc_kernel = 8'h03;
     14'b10010010100010: fc_kernel = 8'h00;
     14'b10010010100011: fc_kernel = 8'hff;
     14'b10010010100100: fc_kernel = 8'hfa;
     14'b10010010100101: fc_kernel = 8'hf0;
     14'b10010010100110: fc_kernel = 8'hed;
     14'b10010010100111: fc_kernel = 8'he1;
     14'b10010010101000: fc_kernel = 8'he1;
     14'b10010010101001: fc_kernel = 8'he3;
     14'b10010010101010: fc_kernel = 8'he7;
     14'b10010010101011: fc_kernel = 8'hf8;
     14'b10010010101100: fc_kernel = 8'hff;
     14'b10010010101101: fc_kernel = 8'h00;
     14'b10010010101110: fc_kernel = 8'hfe;
     14'b10010010101111: fc_kernel = 8'hfe;
     14'b10010010110000: fc_kernel = 8'h05;
     14'b10010010110001: fc_kernel = 8'hfd;
     14'b10010010110010: fc_kernel = 8'h02;
     14'b10010010110011: fc_kernel = 8'h03;
     14'b10010010110100: fc_kernel = 8'h0a;
     14'b10010010110101: fc_kernel = 8'h0a;
     14'b10010010110110: fc_kernel = 8'h00;
     14'b10010010110111: fc_kernel = 8'hff;
     14'b10010010111000: fc_kernel = 8'hfb;
     14'b10010010111001: fc_kernel = 8'hfe;
     14'b10010010111010: fc_kernel = 8'hfc;
     14'b10010010111011: fc_kernel = 8'hfc;
     14'b10010010111100: fc_kernel = 8'hf7;
     14'b10010010111101: fc_kernel = 8'hf8;
     14'b10010010111110: fc_kernel = 8'heb;
     14'b10010010111111: fc_kernel = 8'he2;
     14'b10010011000000: fc_kernel = 8'he7;
     14'b10010011000001: fc_kernel = 8'hea;
     14'b10010011000010: fc_kernel = 8'hee;
     14'b10010011000011: fc_kernel = 8'h01;
     14'b10010011000100: fc_kernel = 8'h01;
     14'b10010011000101: fc_kernel = 8'h06;
     14'b10010011000110: fc_kernel = 8'h00;
     14'b10010011000111: fc_kernel = 8'h00;
     14'b10010011001000: fc_kernel = 8'h01;
     14'b10010011001001: fc_kernel = 8'h02;
     14'b10010011001010: fc_kernel = 8'h07;
     14'b10010011001011: fc_kernel = 8'h01;
     14'b10010011001100: fc_kernel = 8'h01;
     14'b10010011001101: fc_kernel = 8'h00;
     14'b10010011001110: fc_kernel = 8'hfc;
     14'b10010011001111: fc_kernel = 8'h01;
     14'b10010011010000: fc_kernel = 8'h04;
     14'b10010011010001: fc_kernel = 8'hff;
     14'b10010011010010: fc_kernel = 8'hfd;
     14'b10010011010011: fc_kernel = 8'hf9;
     14'b10010011010100: fc_kernel = 8'hf7;
     14'b10010011010101: fc_kernel = 8'hee;
     14'b10010011010110: fc_kernel = 8'heb;
     14'b10010011010111: fc_kernel = 8'he3;
     14'b10010011011000: fc_kernel = 8'hdd;
     14'b10010011011001: fc_kernel = 8'he7;
     14'b10010011011010: fc_kernel = 8'hfd;
     14'b10010011011011: fc_kernel = 8'h00;
     14'b10010011011100: fc_kernel = 8'h09;
     14'b10010011011101: fc_kernel = 8'h04;
     14'b10010011011110: fc_kernel = 8'h05;
     14'b10010011011111: fc_kernel = 8'h0a;
     14'b10010011100000: fc_kernel = 8'h09;
     14'b10010011100001: fc_kernel = 8'h10;
     14'b10010011100010: fc_kernel = 8'h0b;
     14'b10010011100011: fc_kernel = 8'h05;
     14'b10010011100100: fc_kernel = 8'h04;
     14'b10010011100101: fc_kernel = 8'h01;
     14'b10010011100110: fc_kernel = 8'h06;
     14'b10010011100111: fc_kernel = 8'h0a;
     14'b10010011101000: fc_kernel = 8'h06;
     14'b10010011101001: fc_kernel = 8'h06;
     14'b10010011101010: fc_kernel = 8'h06;
     14'b10010011101011: fc_kernel = 8'h05;
     14'b10010011101100: fc_kernel = 8'hf9;
     14'b10010011101101: fc_kernel = 8'hf6;
     14'b10010011101110: fc_kernel = 8'he2;
     14'b10010011101111: fc_kernel = 8'hdc;
     14'b10010011110000: fc_kernel = 8'hdb;
     14'b10010011110001: fc_kernel = 8'hf5;
     14'b10010011110010: fc_kernel = 8'h0a;
     14'b10010011110011: fc_kernel = 8'h07;
     14'b10010011110100: fc_kernel = 8'h05;
     14'b10010011110101: fc_kernel = 8'h0b;
     14'b10010011110110: fc_kernel = 8'h07;
     14'b10010011110111: fc_kernel = 8'h0c;
     14'b10010011111000: fc_kernel = 8'h08;
     14'b10010011111001: fc_kernel = 8'h07;
     14'b10010011111010: fc_kernel = 8'hf9;
     14'b10010011111011: fc_kernel = 8'h00;
     14'b10010011111100: fc_kernel = 8'h07;
     14'b10010011111101: fc_kernel = 8'h08;
     14'b10010011111110: fc_kernel = 8'h0e;
     14'b10010011111111: fc_kernel = 8'h0f;
     14'b10010100000000: fc_kernel = 8'h0a;
     14'b10010100000001: fc_kernel = 8'h0b;
     14'b10010100000010: fc_kernel = 8'h12;
     14'b10010100000011: fc_kernel = 8'h0e;
     14'b10010100000100: fc_kernel = 8'h0d;
     14'b10010100000101: fc_kernel = 8'h03;
     14'b10010100000110: fc_kernel = 8'he8;
     14'b10010100000111: fc_kernel = 8'hbd;
     14'b10010100001000: fc_kernel = 8'he5;
     14'b10010100001001: fc_kernel = 8'hfe;
     14'b10010100001010: fc_kernel = 8'h0f;
     14'b10010100001011: fc_kernel = 8'h0f;
     14'b10010100001100: fc_kernel = 8'h0d;
     14'b10010100001101: fc_kernel = 8'h07;
     14'b10010100001110: fc_kernel = 8'h07;
     14'b10010100001111: fc_kernel = 8'h05;
     14'b10010100010000: fc_kernel = 8'h07;
     14'b10010100010001: fc_kernel = 8'hff;
     14'b10010100010010: fc_kernel = 8'hf4;
     14'b10010100010011: fc_kernel = 8'h03;
     14'b10010100010100: fc_kernel = 8'h09;
     14'b10010100010101: fc_kernel = 8'h0d;
     14'b10010100010110: fc_kernel = 8'h10;
     14'b10010100010111: fc_kernel = 8'h09;
     14'b10010100011000: fc_kernel = 8'h0d;
     14'b10010100011001: fc_kernel = 8'h0b;
     14'b10010100011010: fc_kernel = 8'h0f;
     14'b10010100011011: fc_kernel = 8'h08;
     14'b10010100011100: fc_kernel = 8'h09;
     14'b10010100011101: fc_kernel = 8'hfb;
     14'b10010100011110: fc_kernel = 8'he4;
     14'b10010100011111: fc_kernel = 8'hb5;
     14'b10010100100000: fc_kernel = 8'hf3;
     14'b10010100100001: fc_kernel = 8'h08;
     14'b10010100100010: fc_kernel = 8'h09;
     14'b10010100100011: fc_kernel = 8'h0b;
     14'b10010100100100: fc_kernel = 8'h07;
     14'b10010100100101: fc_kernel = 8'h09;
     14'b10010100100110: fc_kernel = 8'h06;
     14'b10010100100111: fc_kernel = 8'h03;
     14'b10010100101000: fc_kernel = 8'h03;
     14'b10010100101001: fc_kernel = 8'hfe;
     14'b10010100101010: fc_kernel = 8'hfb;
     14'b10010100101011: fc_kernel = 8'h05;
     14'b10010100101100: fc_kernel = 8'h01;
     14'b10010100101101: fc_kernel = 8'h06;
     14'b10010100101110: fc_kernel = 8'h0d;
     14'b10010100101111: fc_kernel = 8'h0a;
     14'b10010100110000: fc_kernel = 8'h04;
     14'b10010100110001: fc_kernel = 8'h0a;
     14'b10010100110010: fc_kernel = 8'h0c;
     14'b10010100110011: fc_kernel = 8'h0a;
     14'b10010100110100: fc_kernel = 8'hff;
     14'b10010100110101: fc_kernel = 8'he9;
     14'b10010100110110: fc_kernel = 8'hcf;
     14'b10010100110111: fc_kernel = 8'hb5;
     14'b10010100111000: fc_kernel = 8'hfd;
     14'b10010100111001: fc_kernel = 8'h0a;
     14'b10010100111010: fc_kernel = 8'h06;
     14'b10010100111011: fc_kernel = 8'h04;
     14'b10010100111100: fc_kernel = 8'h08;
     14'b10010100111101: fc_kernel = 8'h02;
     14'b10010100111110: fc_kernel = 8'h03;
     14'b10010100111111: fc_kernel = 8'hfe;
     14'b10010101000000: fc_kernel = 8'hfe;
     14'b10010101000001: fc_kernel = 8'hfe;
     14'b10010101000010: fc_kernel = 8'h00;
     14'b10010101000011: fc_kernel = 8'hfb;
     14'b10010101000100: fc_kernel = 8'hf8;
     14'b10010101000101: fc_kernel = 8'h09;
     14'b10010101000110: fc_kernel = 8'h0b;
     14'b10010101000111: fc_kernel = 8'h0c;
     14'b10010101001000: fc_kernel = 8'h02;
     14'b10010101001001: fc_kernel = 8'hff;
     14'b10010101001010: fc_kernel = 8'h05;
     14'b10010101001011: fc_kernel = 8'h03;
     14'b10010101001100: fc_kernel = 8'hfe;
     14'b10010101001101: fc_kernel = 8'he8;
     14'b10010101001110: fc_kernel = 8'hc5;
     14'b10010101001111: fc_kernel = 8'hb0;
     14'b10010101010000: fc_kernel = 8'hfa;
     14'b10010101010001: fc_kernel = 8'h04;
     14'b10010101010010: fc_kernel = 8'h02;
     14'b10010101010011: fc_kernel = 8'hfe;
     14'b10010101010100: fc_kernel = 8'h02;
     14'b10010101010101: fc_kernel = 8'h02;
     14'b10010101010110: fc_kernel = 8'h02;
     14'b10010101010111: fc_kernel = 8'hfd;
     14'b10010101011000: fc_kernel = 8'hfd;
     14'b10010101011001: fc_kernel = 8'h02;
     14'b10010101011010: fc_kernel = 8'hff;
     14'b10010101011011: fc_kernel = 8'hf6;
     14'b10010101011100: fc_kernel = 8'hfe;
     14'b10010101011101: fc_kernel = 8'h02;
     14'b10010101011110: fc_kernel = 8'h0a;
     14'b10010101011111: fc_kernel = 8'h06;
     14'b10010101100000: fc_kernel = 8'h03;
     14'b10010101100001: fc_kernel = 8'hfb;
     14'b10010101100010: fc_kernel = 8'hf7;
     14'b10010101100011: fc_kernel = 8'hf5;
     14'b10010101100100: fc_kernel = 8'hf4;
     14'b10010101100101: fc_kernel = 8'hec;
     14'b10010101100110: fc_kernel = 8'hcf;
     14'b10010101100111: fc_kernel = 8'hb2;
     14'b10010101101000: fc_kernel = 8'he3;
     14'b10010101101001: fc_kernel = 8'hf3;
     14'b10010101101010: fc_kernel = 8'hfd;
     14'b10010101101011: fc_kernel = 8'hfa;
     14'b10010101101100: fc_kernel = 8'hf7;
     14'b10010101101101: fc_kernel = 8'h02;
     14'b10010101101110: fc_kernel = 8'h02;
     14'b10010101101111: fc_kernel = 8'hfc;
     14'b10010101110000: fc_kernel = 8'h02;
     14'b10010101110001: fc_kernel = 8'h00;
     14'b10010101110010: fc_kernel = 8'hfc;
     14'b10010101110011: fc_kernel = 8'hf4;
     14'b10010101110100: fc_kernel = 8'h00;
     14'b10010101110101: fc_kernel = 8'h02;
     14'b10010101110110: fc_kernel = 8'h04;
     14'b10010101110111: fc_kernel = 8'h07;
     14'b10010101111000: fc_kernel = 8'h01;
     14'b10010101111001: fc_kernel = 8'hfa;
     14'b10010101111010: fc_kernel = 8'hf5;
     14'b10010101111011: fc_kernel = 8'hf8;
     14'b10010101111100: fc_kernel = 8'hf7;
     14'b10010101111101: fc_kernel = 8'he5;
     14'b10010101111110: fc_kernel = 8'hd1;
     14'b10010101111111: fc_kernel = 8'hbf;
     14'b10010110000000: fc_kernel = 8'hec;
     14'b10010110000001: fc_kernel = 8'hed;
     14'b10010110000010: fc_kernel = 8'hec;
     14'b10010110000011: fc_kernel = 8'heb;
     14'b10010110000100: fc_kernel = 8'hf6;
     14'b10010110000101: fc_kernel = 8'hff;
     14'b10010110000110: fc_kernel = 8'h00;
     14'b10010110000111: fc_kernel = 8'h00;
     14'b10010110001000: fc_kernel = 8'h04;
     14'b10010110001001: fc_kernel = 8'h04;
     14'b10010110001010: fc_kernel = 8'hf4;
     14'b10010110001011: fc_kernel = 8'hf6;
     14'b10010110001100: fc_kernel = 8'hff;
     14'b10010110001101: fc_kernel = 8'h06;
     14'b10010110001110: fc_kernel = 8'h02;
     14'b10010110001111: fc_kernel = 8'h02;
     14'b10010110010000: fc_kernel = 8'hfc;
     14'b10010110010001: fc_kernel = 8'h00;
     14'b10010110010010: fc_kernel = 8'hfc;
     14'b10010110010011: fc_kernel = 8'hf8;
     14'b10010110010100: fc_kernel = 8'hed;
     14'b10010110010101: fc_kernel = 8'he0;
     14'b10010110010110: fc_kernel = 8'hca;
     14'b10010110010111: fc_kernel = 8'hc4;
     14'b10010110011000: fc_kernel = 8'he4;
     14'b10010110011001: fc_kernel = 8'hdf;
     14'b10010110011010: fc_kernel = 8'hec;
     14'b10010110011011: fc_kernel = 8'hef;
     14'b10010110011100: fc_kernel = 8'hfb;
     14'b10010110011101: fc_kernel = 8'hfd;
     14'b10010110011110: fc_kernel = 8'hf3;
     14'b10010110011111: fc_kernel = 8'hf5;
     14'b10010110100000: fc_kernel = 8'hf9;
     14'b10010110100001: fc_kernel = 8'hfa;
     14'b10010110100010: fc_kernel = 8'hf1;
     14'b10010110100011: fc_kernel = 8'hf8;
     14'b10010110100100: fc_kernel = 8'hfb;
     14'b10010110100101: fc_kernel = 8'h00;
     14'b10010110100110: fc_kernel = 8'hfe;
     14'b10010110100111: fc_kernel = 8'hfc;
     14'b10010110101000: fc_kernel = 8'hf5;
     14'b10010110101001: fc_kernel = 8'hfd;
     14'b10010110101010: fc_kernel = 8'hf9;
     14'b10010110101011: fc_kernel = 8'hf5;
     14'b10010110101100: fc_kernel = 8'hed;
     14'b10010110101101: fc_kernel = 8'he7;
     14'b10010110101110: fc_kernel = 8'he6;
     14'b10010110101111: fc_kernel = 8'hde;
     14'b10010110110000: fc_kernel = 8'hd1;
     14'b10010110110001: fc_kernel = 8'hdf;
     14'b10010110110010: fc_kernel = 8'hf3;
     14'b10010110110011: fc_kernel = 8'hfb;
     14'b10010110110100: fc_kernel = 8'hfd;
     14'b10010110110101: fc_kernel = 8'hf6;
     14'b10010110110110: fc_kernel = 8'hf4;
     14'b10010110110111: fc_kernel = 8'hef;
     14'b10010110111000: fc_kernel = 8'heb;
     14'b10010110111001: fc_kernel = 8'he5;
     14'b10010110111010: fc_kernel = 8'hea;
     14'b10010110111011: fc_kernel = 8'hf2;
     14'b10010110111100: fc_kernel = 8'hfa;
     14'b10010110111101: fc_kernel = 8'hf9;
     14'b10010110111110: fc_kernel = 8'hfb;
     14'b10010110111111: fc_kernel = 8'hf6;
     14'b10010111000000: fc_kernel = 8'hf9;
     14'b10010111000001: fc_kernel = 8'hfd;
     14'b10010111000010: fc_kernel = 8'hfb;
     14'b10010111000011: fc_kernel = 8'hf2;
     14'b10010111000100: fc_kernel = 8'he3;
     14'b10010111000101: fc_kernel = 8'hea;
     14'b10010111000110: fc_kernel = 8'hf7;
     14'b10010111000111: fc_kernel = 8'hfc;
     14'b10010111001000: fc_kernel = 8'hd4;
     14'b10010111001001: fc_kernel = 8'hea;
     14'b10010111001010: fc_kernel = 8'hff;
     14'b10010111001011: fc_kernel = 8'h04;
     14'b10010111001100: fc_kernel = 8'h00;
     14'b10010111001101: fc_kernel = 8'hfb;
     14'b10010111001110: fc_kernel = 8'hf8;
     14'b10010111001111: fc_kernel = 8'hf6;
     14'b10010111010000: fc_kernel = 8'hf2;
     14'b10010111010001: fc_kernel = 8'hed;
     14'b10010111010010: fc_kernel = 8'hec;
     14'b10010111010011: fc_kernel = 8'hf5;
     14'b10010111010100: fc_kernel = 8'hf3;
     14'b10010111010101: fc_kernel = 8'hf7;
     14'b10010111010110: fc_kernel = 8'hfa;
     14'b10010111010111: fc_kernel = 8'hf5;
     14'b10010111011000: fc_kernel = 8'hf2;
     14'b10010111011001: fc_kernel = 8'hf4;
     14'b10010111011010: fc_kernel = 8'hf8;
     14'b10010111011011: fc_kernel = 8'hee;
     14'b10010111011100: fc_kernel = 8'he3;
     14'b10010111011101: fc_kernel = 8'hf1;
     14'b10010111011110: fc_kernel = 8'hfe;
     14'b10010111011111: fc_kernel = 8'h05;
     14'b10010111100000: fc_kernel = 8'hf8;
     14'b10010111100001: fc_kernel = 8'h00;
     14'b10010111100010: fc_kernel = 8'hf9;
     14'b10010111100011: fc_kernel = 8'hf9;
     14'b10010111100100: fc_kernel = 8'hf2;
     14'b10010111100101: fc_kernel = 8'hf5;
     14'b10010111100110: fc_kernel = 8'hf7;
     14'b10010111100111: fc_kernel = 8'hfc;
     14'b10010111101000: fc_kernel = 8'hfa;
     14'b10010111101001: fc_kernel = 8'hf9;
     14'b10010111101010: fc_kernel = 8'hfb;
     14'b10010111101011: fc_kernel = 8'hf8;
     14'b10010111101100: fc_kernel = 8'hfa;
     14'b10010111101101: fc_kernel = 8'hf7;
     14'b10010111101110: fc_kernel = 8'hfb;
     14'b10010111101111: fc_kernel = 8'hf3;
     14'b10010111110000: fc_kernel = 8'hf0;
     14'b10010111110001: fc_kernel = 8'hf2;
     14'b10010111110010: fc_kernel = 8'hef;
     14'b10010111110011: fc_kernel = 8'hf6;
     14'b10010111110100: fc_kernel = 8'hf0;
     14'b10010111110101: fc_kernel = 8'hfb;
     14'b10010111110110: fc_kernel = 8'h05;
     14'b10010111110111: fc_kernel = 8'h0a;
     14'b10010111111000: fc_kernel = 8'hf0;
     14'b10010111111001: fc_kernel = 8'h00;
     14'b10010111111010: fc_kernel = 8'hf4;
     14'b10010111111011: fc_kernel = 8'hec;
     14'b10010111111100: fc_kernel = 8'heb;
     14'b10010111111101: fc_kernel = 8'hf6;
     14'b10010111111110: fc_kernel = 8'hf6;
     14'b10010111111111: fc_kernel = 8'hf5;
     14'b10011000000000: fc_kernel = 8'hf2;
     14'b10011000000001: fc_kernel = 8'hf9;
     14'b10011000000010: fc_kernel = 8'hf2;
     14'b10011000000011: fc_kernel = 8'hf7;
     14'b10011000000100: fc_kernel = 8'hf5;
     14'b10011000000101: fc_kernel = 8'hf7;
     14'b10011000000110: fc_kernel = 8'hf0;
     14'b10011000000111: fc_kernel = 8'hf7;
     14'b10011000001000: fc_kernel = 8'hf3;
     14'b10011000001001: fc_kernel = 8'hf4;
     14'b10011000001010: fc_kernel = 8'hf3;
     14'b10011000001011: fc_kernel = 8'hf7;
     14'b10011000001100: fc_kernel = 8'hfe;
     14'b10011000001101: fc_kernel = 8'h0c;
     14'b10011000001110: fc_kernel = 8'h08;
     14'b10011000001111: fc_kernel = 8'h08;
     14'b10011000010000: fc_kernel = 8'hfc;
     14'b10011000010001: fc_kernel = 8'hfa;
     14'b10011000010010: fc_kernel = 8'hff;
     14'b10011000010011: fc_kernel = 8'hff;
     14'b10011000010100: fc_kernel = 8'hfa;
     14'b10011000010101: fc_kernel = 8'h00;
     14'b10011000010110: fc_kernel = 8'h01;
     14'b10011000010111: fc_kernel = 8'hfd;
     14'b10011000011000: fc_kernel = 8'hfe;
     14'b10011000011001: fc_kernel = 8'hfa;
     14'b10011000011010: fc_kernel = 8'hfa;
     14'b10011000011011: fc_kernel = 8'hf3;
     14'b10011000011100: fc_kernel = 8'hf3;
     14'b10011000011101: fc_kernel = 8'hf8;
     14'b10011000011110: fc_kernel = 8'hfd;
     14'b10011000011111: fc_kernel = 8'hfe;
     14'b10011000100000: fc_kernel = 8'hf8;
     14'b10011000100001: fc_kernel = 8'hfd;
     14'b10011000100010: fc_kernel = 8'h05;
     14'b10011000100011: fc_kernel = 8'h0a;
     14'b10011000100100: fc_kernel = 8'h08;
     14'b10011000100101: fc_kernel = 8'h0c;
     14'b10011000100110: fc_kernel = 8'h01;
     14'b10011000100111: fc_kernel = 8'hf1;
     14'b10011000101000: fc_kernel = 8'hf6;
     14'b10011000101001: fc_kernel = 8'hf9;
     14'b10011000101010: fc_kernel = 8'h0e;
     14'b10011000101011: fc_kernel = 8'h19;
     14'b10011000101100: fc_kernel = 8'h21;
     14'b10011000101101: fc_kernel = 8'h18;
     14'b10011000101110: fc_kernel = 8'h15;
     14'b10011000101111: fc_kernel = 8'h11;
     14'b10011000110000: fc_kernel = 8'h0e;
     14'b10011000110001: fc_kernel = 8'h0f;
     14'b10011000110010: fc_kernel = 8'h0e;
     14'b10011000110011: fc_kernel = 8'h0c;
     14'b10011000110100: fc_kernel = 8'h0c;
     14'b10011000110101: fc_kernel = 8'h0c;
     14'b10011000110110: fc_kernel = 8'h0d;
     14'b10011000110111: fc_kernel = 8'h10;
     14'b10011000111000: fc_kernel = 8'h0c;
     14'b10011000111001: fc_kernel = 8'h14;
     14'b10011000111010: fc_kernel = 8'h1a;
     14'b10011000111011: fc_kernel = 8'h19;
     14'b10011000111100: fc_kernel = 8'h10;
     14'b10011000111101: fc_kernel = 8'h06;
     14'b10011000111110: fc_kernel = 8'h00;
     14'b10011000111111: fc_kernel = 8'hf3;
     default: fc_kernel = 8'h0;
    endcase
    end

endfunction